* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lcesd1_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT lcesd2_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_shield PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_wos PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_x_40k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_x_40k PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_x_40k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nr36 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_w40 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pad_corner
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_70
** N=4 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT padbox
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pad_in VSS pad VDD DataIn
** N=24 EP=4 IP=1 FDC=96
M0 VSS VSS 7 VSS N L=3.5e-07 W=9e-06 $X=5700 $Y=147100 $D=0
M1 8 7 VSS VSS N L=3.5e-07 W=9e-06 $X=8100 $Y=147100 $D=0
M2 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=13200 $Y=147100 $D=0
M3 10 VSS VSS VSS N L=3.5e-07 W=9e-06 $X=15600 $Y=147100 $D=0
M4 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=191300 $D=0
M5 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=196210 $D=0
M6 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=197780 $D=0
M7 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=202690 $D=0
M8 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=204260 $D=0
M9 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=209170 $D=0
M10 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=210740 $D=0
M11 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=215650 $D=0
M12 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=217220 $D=0
M13 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=222130 $D=0
M14 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=18000 $Y=147100 $D=0
M15 10 VSS VSS VSS N L=3.5e-07 W=9e-06 $X=20400 $Y=147100 $D=0
M16 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=22800 $Y=147100 $D=0
M17 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=25200 $Y=147100 $D=0
M18 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=27600 $Y=147100 $D=0
M19 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=30000 $Y=147100 $D=0
M20 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=32400 $Y=147100 $D=0
M21 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=34800 $Y=147100 $D=0
M22 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=37200 $Y=147100 $D=0
M23 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=39600 $Y=147100 $D=0
M24 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=42000 $Y=147100 $D=0
M25 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=44400 $Y=147100 $D=0
M26 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=191300 $D=0
M27 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=196210 $D=0
M28 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=197780 $D=0
M29 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=202690 $D=0
M30 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=204260 $D=0
M31 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=209170 $D=0
M32 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=210740 $D=0
M33 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=215650 $D=0
M34 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=217220 $D=0
M35 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=222130 $D=0
M36 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=59400 $Y=146950 $D=0
M37 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=61800 $Y=146950 $D=0
M38 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=64200 $Y=146950 $D=0
M39 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=66600 $Y=146950 $D=0
M40 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=69000 $Y=146950 $D=0
M41 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=71400 $Y=146950 $D=0
M42 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=73800 $Y=146950 $D=0
M43 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=76200 $Y=146950 $D=0
M44 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=78600 $Y=146950 $D=0
M45 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=81000 $Y=146950 $D=0
M46 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=83400 $Y=146950 $D=0
M47 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=85800 $Y=146950 $D=0
M48 VDD VSS 7 VDD P L=3.5e-07 W=1.56e-05 $X=5700 $Y=165550 $D=16
M49 8 7 VDD VDD P L=3.5e-07 W=1.56e-05 $X=8100 $Y=165550 $D=16
M50 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=13200 $Y=165550 $D=16
M51 9 VSS VDD VDD P L=3.5e-07 W=1.56e-05 $X=15600 $Y=165550 $D=16
M52 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=97085 $D=16
M53 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=101995 $D=16
M54 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=103565 $D=16
M55 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=108475 $D=16
M56 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=110045 $D=16
M57 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=114955 $D=16
M58 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=116525 $D=16
M59 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=121435 $D=16
M60 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=123005 $D=16
M61 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=127915 $D=16
M62 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=18000 $Y=165550 $D=16
M63 9 VSS VDD VDD P L=3.5e-07 W=1.56e-05 $X=20400 $Y=165550 $D=16
M64 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=22800 $Y=165550 $D=16
M65 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=25200 $Y=165550 $D=16
M66 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=27600 $Y=165550 $D=16
M67 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=30000 $Y=165550 $D=16
M68 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=32400 $Y=165550 $D=16
M69 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=34800 $Y=165550 $D=16
M70 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=37200 $Y=165550 $D=16
M71 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=39600 $Y=165550 $D=16
M72 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=42000 $Y=165550 $D=16
M73 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=44400 $Y=165550 $D=16
M74 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=97085 $D=16
M75 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=101995 $D=16
M76 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=103565 $D=16
M77 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=108475 $D=16
M78 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=110045 $D=16
M79 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=114955 $D=16
M80 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=116525 $D=16
M81 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=121435 $D=16
M82 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=123005 $D=16
M83 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=127915 $D=16
M84 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=59400 $Y=165550 $D=16
M85 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=61800 $Y=165550 $D=16
M86 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=64200 $Y=165550 $D=16
M87 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=66600 $Y=165550 $D=16
M88 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=69000 $Y=165550 $D=16
M89 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=71400 $Y=165550 $D=16
M90 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=73800 $Y=165550 $D=16
M91 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=76200 $Y=165550 $D=16
M92 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=78600 $Y=165550 $D=16
M93 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=81000 $Y=165550 $D=16
M94 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=83400 $Y=165550 $D=16
M95 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=85800 $Y=165550 $D=16
.ENDS
***************************************
.SUBCKT pad_out VDD DataOut pad VSS
** N=25 EP=4 IP=1 FDC=96
M0 VSS VDD 7 VSS N L=3.5e-07 W=9e-06 $X=5700 $Y=147100 $D=0
M1 8 7 VSS VSS N L=3.5e-07 W=9e-06 $X=8100 $Y=147100 $D=0
M2 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=13200 $Y=147100 $D=0
M3 10 DataOut VSS VSS N L=3.5e-07 W=9e-06 $X=15600 $Y=147100 $D=0
M4 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=191300 $D=0
M5 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=196210 $D=0
M6 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=197780 $D=0
M7 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=202690 $D=0
M8 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=204260 $D=0
M9 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=209170 $D=0
M10 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=210740 $D=0
M11 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=215650 $D=0
M12 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=217220 $D=0
M13 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=222130 $D=0
M14 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=18000 $Y=147100 $D=0
M15 10 DataOut VSS VSS N L=3.5e-07 W=9e-06 $X=20400 $Y=147100 $D=0
M16 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=22800 $Y=147100 $D=0
M17 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=25200 $Y=147100 $D=0
M18 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=27600 $Y=147100 $D=0
M19 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=30000 $Y=147100 $D=0
M20 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=32400 $Y=147100 $D=0
M21 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=34800 $Y=147100 $D=0
M22 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=37200 $Y=147100 $D=0
M23 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=39600 $Y=147100 $D=0
M24 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=42000 $Y=147100 $D=0
M25 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=44400 $Y=147100 $D=0
M26 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=191300 $D=0
M27 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=196210 $D=0
M28 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=197780 $D=0
M29 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=202690 $D=0
M30 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=204260 $D=0
M31 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=209170 $D=0
M32 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=210740 $D=0
M33 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=215650 $D=0
M34 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=217220 $D=0
M35 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=222130 $D=0
M36 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=59400 $Y=146950 $D=0
M37 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=61800 $Y=146950 $D=0
M38 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=64200 $Y=146950 $D=0
M39 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=66600 $Y=146950 $D=0
M40 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=69000 $Y=146950 $D=0
M41 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=71400 $Y=146950 $D=0
M42 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=73800 $Y=146950 $D=0
M43 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=76200 $Y=146950 $D=0
M44 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=78600 $Y=146950 $D=0
M45 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=81000 $Y=146950 $D=0
M46 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=83400 $Y=146950 $D=0
M47 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=85800 $Y=146950 $D=0
M48 VDD VDD 7 VDD P L=3.5e-07 W=1.56e-05 $X=5700 $Y=165550 $D=16
M49 8 7 VDD VDD P L=3.5e-07 W=1.56e-05 $X=8100 $Y=165550 $D=16
M50 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=13200 $Y=165550 $D=16
M51 9 DataOut VDD VDD P L=3.5e-07 W=1.56e-05 $X=15600 $Y=165550 $D=16
M52 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=97085 $D=16
M53 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=101995 $D=16
M54 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=103565 $D=16
M55 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=108475 $D=16
M56 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=110045 $D=16
M57 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=114955 $D=16
M58 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=116525 $D=16
M59 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=121435 $D=16
M60 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=123005 $D=16
M61 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=127915 $D=16
M62 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=18000 $Y=165550 $D=16
M63 9 DataOut VDD VDD P L=3.5e-07 W=1.56e-05 $X=20400 $Y=165550 $D=16
M64 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=22800 $Y=165550 $D=16
M65 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=25200 $Y=165550 $D=16
M66 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=27600 $Y=165550 $D=16
M67 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=30000 $Y=165550 $D=16
M68 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=32400 $Y=165550 $D=16
M69 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=34800 $Y=165550 $D=16
M70 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=37200 $Y=165550 $D=16
M71 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=39600 $Y=165550 $D=16
M72 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=42000 $Y=165550 $D=16
M73 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=44400 $Y=165550 $D=16
M74 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=97085 $D=16
M75 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=101995 $D=16
M76 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=103565 $D=16
M77 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=108475 $D=16
M78 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=110045 $D=16
M79 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=114955 $D=16
M80 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=116525 $D=16
M81 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=121435 $D=16
M82 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=123005 $D=16
M83 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=127915 $D=16
M84 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=59400 $Y=165550 $D=16
M85 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=61800 $Y=165550 $D=16
M86 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=64200 $Y=165550 $D=16
M87 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=66600 $Y=165550 $D=16
M88 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=69000 $Y=165550 $D=16
M89 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=71400 $Y=165550 $D=16
M90 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=73800 $Y=165550 $D=16
M91 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=76200 $Y=165550 $D=16
M92 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=78600 $Y=165550 $D=16
M93 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=81000 $Y=165550 $D=16
M94 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=83400 $Y=165550 $D=16
M95 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=85800 $Y=165550 $D=16
.ENDS
***************************************
.SUBCKT ICV_69 1 2 3 4 5
** N=7 EP=5 IP=12 FDC=192
X0 1 4 2 3 pad_in $T=0 323200 0 270 $X=0 $Y=232300
X1 2 1 5 1 pad_out $T=0 413200 0 270 $X=0 $Y=322300
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 5
** N=7 EP=4 IP=6 FDC=96
X0 2 3 5 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_68
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1 VSS VDD
** N=38 EP=2 IP=1 FDC=1
D0 VSS VDD pdio_m AREA=9e-10 PJ=0.00012 $X=8570 $Y=96300 $D=31
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3
** N=5 EP=3 IP=6 FDC=96
X0 2 1 3 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_67 1 2 3 4
** N=6 EP=4 IP=12 FDC=192
X0 2 1 3 1 pad_out $T=0 773200 0 270 $X=0 $Y=682300
X1 2 1 4 1 pad_out $T=0 863200 0 270 $X=0 $Y=772300
.ENDS
***************************************
.SUBCKT ICV_66 1 2 3 4
** N=6 EP=4 IP=12 FDC=192
X0 2 1 3 1 pad_out $T=0 953200 0 270 $X=0 $Y=862300
X1 2 1 4 1 pad_out $T=0 1043200 0 270 $X=0 $Y=952300
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3
** N=5 EP=3 IP=6 FDC=96
X0 2 1 3 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_65 1 2 3 4
** N=6 EP=4 IP=12 FDC=192
X0 2 1 3 1 pad_out $T=0 1223200 0 270 $X=0 $Y=1132300
X1 2 1 4 1 pad_out $T=0 1313200 0 270 $X=0 $Y=1222300
.ENDS
***************************************
.SUBCKT ICV_64 1 2 3
** N=5 EP=3 IP=10 FDC=96
X1 2 1 3 1 pad_out $T=0 1403200 0 270 $X=0 $Y=1312300
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
** N=21 EP=19 IP=88 FDC=1344
X1 1 6 2 3 pad_in $T=323200 1636400 0 180 $X=232300 $Y=1402300
X2 2 1 7 1 pad_out $T=503200 1636400 0 180 $X=412300 $Y=1402300
X3 2 1 8 1 pad_out $T=593200 1636400 0 180 $X=502300 $Y=1402300
X4 2 1 9 1 pad_out $T=683200 1636400 0 180 $X=592300 $Y=1402300
X5 2 4 10 1 pad_out $T=773200 1636400 0 180 $X=682300 $Y=1402300
X6 2 1 11 1 pad_out $T=863200 1636400 0 180 $X=772300 $Y=1402300
X7 2 5 12 1 pad_out $T=953200 1636400 0 180 $X=862300 $Y=1402300
X8 2 1 13 1 pad_out $T=1043200 1636400 0 180 $X=952300 $Y=1402300
X9 2 1 14 1 pad_out $T=1133200 1636400 0 180 $X=1042300 $Y=1402300
X10 2 1 15 1 pad_out $T=1223200 1636400 0 180 $X=1132300 $Y=1402300
X11 2 1 16 1 pad_out $T=1313200 1636400 0 180 $X=1222300 $Y=1402300
X12 2 1 17 1 pad_out $T=1403200 1636400 0 180 $X=1312300 $Y=1402300
X13 2 1 18 1 pad_out $T=1493200 1636400 0 180 $X=1402300 $Y=1402300
X14 2 1 19 1 pad_out $T=1726400 1313200 0 90 $X=1492300 $Y=1312300
.ENDS
***************************************
.SUBCKT pad_fill_4
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_01
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_62
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT pad_fill_005
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_60
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_61
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_63 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
** N=21 EP=19 IP=418 FDC=1248
X1 1 7 2 3 pad_in $T=239630 0 0 0 $X=238730 $Y=0
X2 1 8 2 4 pad_in $T=336060 0 0 0 $X=335160 $Y=0
X3 1 9 2 5 pad_in $T=1011050 0 0 0 $X=1010150 $Y=0
X4 2 1 10 1 pad_out $T=432490 0 0 0 $X=431590 $Y=0
X5 2 1 11 1 pad_out $T=528920 0 0 0 $X=528020 $Y=0
X6 2 1 12 1 pad_out $T=625350 0 0 0 $X=624450 $Y=0
X7 2 1 13 1 pad_out $T=721775 0 0 0 $X=720875 $Y=0
X8 2 1 14 1 pad_out $T=818200 0 0 0 $X=817300 $Y=0
X9 2 1 15 1 pad_out $T=914625 0 0 0 $X=913725 $Y=0
X10 2 1 16 1 pad_out $T=1107480 0 0 0 $X=1106580 $Y=0
X11 2 6 17 1 pad_out $T=1203910 0 0 0 $X=1203010 $Y=0
X12 2 1 18 1 pad_out $T=1300340 0 0 0 $X=1299440 $Y=0
X13 2 1 19 1 pad_out $T=1396770 0 0 0 $X=1395870 $Y=0
.ENDS
***************************************
.SUBCKT FILL32
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_44
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_48
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_58
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=5 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT FILL16
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL8
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_52
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT DFFQSRX1 D CLK SETB RESETB VSS VDD Q
** N=34 EP=7 IP=0 FDC=40
M0 VSS D 20 VSS N L=1.8e-07 W=2.2e-07 $X=945 $Y=750 $D=0
M1 10 CLK VSS VSS N L=1.8e-07 W=2.2e-07 $X=1745 $Y=750 $D=0
M2 11 10 20 VSS N L=1.8e-07 W=2.2e-07 $X=3245 $Y=755 $D=0
M3 12 11 VSS VSS N L=1.8e-07 W=2.2e-07 $X=4745 $Y=755 $D=0
M4 13 12 VSS VSS N L=1.8e-07 W=2.2e-07 $X=6250 $Y=760 $D=0
M5 VSS 14 13 VSS N L=1.8e-07 W=2.2e-07 $X=7050 $Y=760 $D=0
M6 15 13 VSS VSS N L=1.8e-07 W=2.2e-07 $X=7850 $Y=1120 $D=0
M7 VSS SETB 14 VSS N L=1.8e-07 W=2.2e-07 $X=9355 $Y=755 $D=0
M8 22 CLK 11 VSS N L=1.8e-07 W=2.2e-07 $X=10860 $Y=750 $D=0
M9 33 15 VSS VSS N L=1.8e-07 W=4.4e-07 $X=12320 $Y=965 $D=0
M10 22 RESETB 33 VSS N L=1.8e-07 W=4.4e-07 $X=13040 $Y=965 $D=0
M11 16 CLK 15 VSS N L=1.8e-07 W=2.2e-07 $X=14500 $Y=755 $D=0
M12 34 16 VSS VSS N L=1.8e-07 W=4.4e-07 $X=15960 $Y=740 $D=0
M13 17 RESETB 34 VSS N L=1.8e-07 W=4.4e-07 $X=16680 $Y=740 $D=0
M14 18 17 VSS VSS N L=1.8e-07 W=2.2e-07 $X=18140 $Y=755 $D=0
M15 19 18 VSS VSS N L=1.8e-07 W=2.2e-07 $X=19640 $Y=755 $D=0
M16 VSS 14 19 VSS N L=1.8e-07 W=2.2e-07 $X=20440 $Y=755 $D=0
M17 24 19 VSS VSS N L=1.8e-07 W=2.2e-07 $X=21240 $Y=755 $D=0
M18 16 10 24 VSS N L=1.8e-07 W=2.2e-07 $X=22740 $Y=755 $D=0
M19 Q 17 VSS VSS N L=1.8e-07 W=2.2e-07 $X=24240 $Y=755 $D=0
M20 VDD D 20 VDD P L=1.8e-07 W=4.4e-07 $X=945 $Y=2705 $D=16
M21 10 CLK VDD VDD P L=1.8e-07 W=4.4e-07 $X=1665 $Y=2705 $D=16
M22 11 CLK 20 VDD P L=1.8e-07 W=4.4e-07 $X=3245 $Y=2725 $D=16
M23 12 11 VDD VDD P L=1.8e-07 W=4.4e-07 $X=4745 $Y=2725 $D=16
M24 21 12 13 VDD P L=1.8e-07 W=8.8e-07 $X=6250 $Y=2300 $D=16
M25 VDD 14 21 VDD P L=1.8e-07 W=8.8e-07 $X=6970 $Y=2300 $D=16
M26 15 13 VDD VDD P L=1.8e-07 W=4.4e-07 $X=7730 $Y=2520 $D=16
M27 VDD SETB 14 VDD P L=1.8e-07 W=4.4e-07 $X=9355 $Y=2535 $D=16
M28 22 10 11 VDD P L=1.8e-07 W=4.4e-07 $X=10815 $Y=2505 $D=16
M29 22 15 VDD VDD P L=1.8e-07 W=4.4e-07 $X=12320 $Y=2505 $D=16
M30 VDD RESETB 22 VDD P L=1.8e-07 W=4.4e-07 $X=13040 $Y=2505 $D=16
M31 16 10 15 VDD P L=1.8e-07 W=4.4e-07 $X=14500 $Y=2505 $D=16
M32 17 16 VDD VDD P L=1.8e-07 W=4.4e-07 $X=15960 $Y=2665 $D=16
M33 VDD RESETB 17 VDD P L=1.8e-07 W=4.4e-07 $X=16680 $Y=2665 $D=16
M34 18 17 VDD VDD P L=1.8e-07 W=4.4e-07 $X=18140 $Y=2725 $D=16
M35 23 18 19 VDD P L=1.8e-07 W=8.8e-07 $X=19640 $Y=2285 $D=16
M36 VDD 14 23 VDD P L=1.8e-07 W=8.8e-07 $X=20360 $Y=2285 $D=16
M37 24 19 VDD VDD P L=1.8e-07 W=4.4e-07 $X=21120 $Y=2505 $D=16
M38 16 CLK 24 VDD P L=1.8e-07 W=4.4e-07 $X=22740 $Y=2505 $D=16
M39 Q 17 VDD VDD P L=1.8e-07 W=4.4e-07 $X=24200 $Y=2505 $D=16
.ENDS
***************************************
.SUBCKT FILL4
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL1
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL2
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT XOR2X1 B A VDD VSS Z
** N=11 EP=5 IP=0 FDC=10
M0 VSS B 10 VSS N L=1.8e-07 W=4.4e-07 $X=630 $Y=985 $D=0
M1 8 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=1350 $Y=985 $D=0
M2 9 8 10 VSS N L=1.8e-07 W=4.4e-07 $X=3205 $Y=1000 $D=0
M3 B A 9 VSS N L=1.8e-07 W=4.4e-07 $X=3925 $Y=1000 $D=0
M4 Z 9 VSS VSS N L=1.8e-07 W=4.4e-07 $X=5345 $Y=1000 $D=0
M5 VDD B 10 VDD P L=1.8e-07 W=4.4e-07 $X=630 $Y=2435 $D=16
M6 8 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1350 $Y=2435 $D=16
M7 9 A 10 VDD P L=1.8e-07 W=4.4e-07 $X=3205 $Y=2435 $D=16
M8 B 8 9 VDD P L=1.8e-07 W=4.4e-07 $X=3925 $Y=2435 $D=16
M9 Z 9 VDD VDD P L=1.8e-07 W=4.4e-07 $X=5345 $Y=2435 $D=16
.ENDS
***************************************
.SUBCKT AND2X1 A B VSS VDD Z
** N=10 EP=5 IP=0 FDC=6
M0 10 A 8 VSS N L=1.8e-07 W=4.4e-07 $X=905 $Y=750 $D=0
M1 VSS B 10 VSS N L=1.8e-07 W=4.4e-07 $X=1625 $Y=750 $D=0
M2 Z 8 VSS VSS N L=1.8e-07 W=2.2e-07 $X=2385 $Y=860 $D=0
M3 8 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=905 $Y=2670 $D=16
M4 VDD B 8 VDD P L=1.8e-07 W=4.4e-07 $X=1625 $Y=2670 $D=16
M5 Z 8 VDD VDD P L=1.8e-07 W=4.4e-07 $X=2385 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT ICV_50
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT OR2X1 A B VSS VDD Z
** N=12 EP=5 IP=0 FDC=6
M0 8 A VSS VSS N L=1.8e-07 W=2.2e-07 $X=835 $Y=760 $D=0
M1 VSS B 8 VSS N L=1.8e-07 W=2.2e-07 $X=1635 $Y=760 $D=0
M2 Z 8 VSS VSS N L=1.8e-07 W=2.2e-07 $X=2435 $Y=760 $D=0
M3 9 A 8 VDD P L=1.8e-07 W=8.8e-07 $X=835 $Y=2300 $D=16
M4 VDD B 9 VDD P L=1.8e-07 W=8.8e-07 $X=1555 $Y=2300 $D=16
M5 Z 8 VDD VDD P L=1.8e-07 W=4.4e-07 $X=2315 $Y=2520 $D=16
.ENDS
***************************************
.SUBCKT NAND3X1 A B C VSS VDD Z
** N=10 EP=6 IP=0 FDC=6
M0 9 A VSS VSS N L=1.8e-07 W=6.6e-07 $X=1210 $Y=745 $D=0
M1 10 B 9 VSS N L=1.8e-07 W=6.6e-07 $X=1930 $Y=745 $D=0
M2 Z C 10 VSS N L=1.8e-07 W=6.6e-07 $X=2650 $Y=745 $D=0
M3 Z A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1210 $Y=2670 $D=16
M4 VDD B Z VDD P L=1.8e-07 W=4.4e-07 $X=1930 $Y=2670 $D=16
M5 Z C VDD VDD P L=1.8e-07 W=4.4e-07 $X=2650 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT NOR2X1 A B VSS VDD Z
** N=10 EP=5 IP=0 FDC=4
M0 Z A VSS VSS N L=1.8e-07 W=2.2e-07 $X=925 $Y=760 $D=0
M1 VSS B Z VSS N L=1.8e-07 W=2.2e-07 $X=1725 $Y=760 $D=0
M2 8 A VDD VDD P L=1.8e-07 W=8.8e-07 $X=925 $Y=2300 $D=16
M3 Z B 8 VDD P L=1.8e-07 W=8.8e-07 $X=1645 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT ICV_37
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT INVX2 A VSS VDD Z
** N=6 EP=4 IP=0 FDC=2
M0 Z A VSS VSS N L=1.8e-07 W=4.4e-07 $X=740 $Y=740 $D=0
M1 Z A VDD VDD P L=1.8e-07 W=8.8e-07 $X=740 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT ICV_51
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT NAND2X1 A B VSS VDD Z
** N=9 EP=5 IP=0 FDC=4
M0 9 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=985 $Y=745 $D=0
M1 Z B 9 VSS N L=1.8e-07 W=4.4e-07 $X=1705 $Y=745 $D=0
M2 Z A VDD VDD P L=1.8e-07 W=4.4e-07 $X=985 $Y=2670 $D=16
M3 VDD B Z VDD P L=1.8e-07 W=4.4e-07 $X=1705 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT ICV_33
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT DFFQX1 CLK Q VDD D VSS
** N=16 EP=5 IP=0 FDC=18
M0 8 CLK VSS VSS N L=1.8e-07 W=2.2e-07 $X=870 $Y=750 $D=0
M1 9 8 D VSS N L=1.8e-07 W=2.2e-07 $X=2370 $Y=750 $D=0
M2 VSS 9 10 VSS N L=1.8e-07 W=2.2e-07 $X=3960 $Y=750 $D=0
M3 12 10 VSS VSS N L=1.8e-07 W=2.2e-07 $X=5720 $Y=750 $D=0
M4 9 CLK 12 VSS N L=1.8e-07 W=2.2e-07 $X=6755 $Y=750 $D=0
M5 11 CLK 10 VSS N L=1.8e-07 W=2.2e-07 $X=8440 $Y=750 $D=0
M6 13 8 11 VSS N L=1.8e-07 W=2.2e-07 $X=9640 $Y=750 $D=0
M7 VSS Q 13 VSS N L=1.8e-07 W=2.2e-07 $X=10440 $Y=750 $D=0
M8 Q 11 VSS VSS N L=1.8e-07 W=2.2e-07 $X=11240 $Y=750 $D=0
M9 8 CLK VDD VDD P L=1.8e-07 W=4.4e-07 $X=870 $Y=2670 $D=16
M10 9 CLK D VDD P L=1.8e-07 W=4.4e-07 $X=2460 $Y=2670 $D=16
M11 VDD 9 10 VDD P L=1.8e-07 W=4.4e-07 $X=3960 $Y=2670 $D=16
M12 12 10 VDD VDD P L=1.8e-07 W=4.4e-07 $X=5460 $Y=2670 $D=16
M13 9 8 12 VDD P L=1.8e-07 W=4.4e-07 $X=6180 $Y=2670 $D=16
M14 11 8 10 VDD P L=1.8e-07 W=4.4e-07 $X=7980 $Y=2670 $D=16
M15 13 CLK 11 VDD P L=1.8e-07 W=4.4e-07 $X=9780 $Y=2670 $D=16
M16 VDD Q 13 VDD P L=1.8e-07 W=4.4e-07 $X=10500 $Y=2670 $D=16
M17 Q 11 VDD VDD P L=1.8e-07 W=4.4e-07 $X=11220 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT ICV_54
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MUX2X1 A S B VSS VDD Z
** N=16 EP=6 IP=0 FDC=12
M0 VSS S 9 VSS N L=1.8e-07 W=4.4e-07 $X=940 $Y=960 $D=0
M1 15 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=1660 $Y=960 $D=0
M2 10 9 15 VSS N L=1.8e-07 W=4.4e-07 $X=2380 $Y=960 $D=0
M3 16 S 10 VSS N L=1.8e-07 W=4.4e-07 $X=3100 $Y=960 $D=0
M4 VSS B 16 VSS N L=1.8e-07 W=4.4e-07 $X=3920 $Y=740 $D=0
M5 Z 10 VSS VSS N L=1.8e-07 W=4.4e-07 $X=4640 $Y=740 $D=0
M6 VDD S 9 VDD P L=1.8e-07 W=4.4e-07 $X=940 $Y=2520 $D=16
M7 11 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1660 $Y=2520 $D=16
M8 10 S 11 VDD P L=1.8e-07 W=4.4e-07 $X=2380 $Y=2520 $D=16
M9 12 9 10 VDD P L=1.8e-07 W=4.4e-07 $X=3100 $Y=2520 $D=16
M10 VDD B 12 VDD P L=1.8e-07 W=4.4e-07 $X=3920 $Y=2735 $D=16
M11 Z 10 VDD VDD P L=1.8e-07 W=4.4e-07 $X=4640 $Y=2735 $D=16
.ENDS
***************************************
.SUBCKT ICV_53
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_56
** N=5 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_59 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
** N=340 EP=37 IP=4747 FDC=3012
X0 1 36 2 268 pad_in $T=1726400 233200 0 90 $X=1492300 $Y=232300
X1 1 37 2 244 pad_in $T=1726400 323200 0 90 $X=1492300 $Y=322300
X249 41 29 34 2 1 2 42 DFFQSRX1 $T=613440 434800 0 0 $X=613010 $Y=434410
X250 48 29 34 2 1 2 46 DFFQSRX1 $T=620160 434800 1 0 $X=619730 $Y=430245
X251 61 29 34 2 1 2 54 DFFQSRX1 $T=667200 434800 1 180 $X=641570 $Y=434410
X252 67 29 34 2 1 2 60 DFFQSRX1 $T=678960 426960 0 180 $X=653330 $Y=422405
X253 74 29 34 2 1 2 62 DFFQSRX1 $T=682880 419120 0 180 $X=657250 $Y=414565
X254 76 29 34 2 1 2 63 DFFQSRX1 $T=682880 458320 0 180 $X=657250 $Y=453765
X255 84 29 34 2 1 2 79 DFFQSRX1 $T=689040 411280 0 0 $X=688610 $Y=410890
X256 97 29 34 2 1 2 86 DFFQSRX1 $T=692400 419120 1 0 $X=691970 $Y=414565
X257 100 29 34 2 1 2 87 DFFQSRX1 $T=722640 426960 1 180 $X=697010 $Y=426570
X258 99 29 34 2 1 2 89 DFFQSRX1 $T=723200 442640 0 180 $X=697570 $Y=438085
X259 101 29 28 2 1 2 106 DFFQSRX1 $T=715360 411280 1 0 $X=714930 $Y=406725
X260 103 29 28 2 1 2 111 DFFQSRX1 $T=715920 403440 1 0 $X=715490 $Y=398885
X261 105 29 28 2 1 2 116 DFFQSRX1 $T=720960 387760 0 0 $X=720530 $Y=387370
X262 127 29 28 2 1 2 130 DFFQSRX1 $T=721520 364240 0 0 $X=721090 $Y=363850
X263 114 29 28 2 1 2 120 DFFQSRX1 $T=721520 372080 0 0 $X=721090 $Y=371690
X264 113 29 28 2 1 2 135 DFFQSRX1 $T=722080 356400 1 0 $X=721650 $Y=351845
X265 109 29 28 2 1 2 121 DFFQSRX1 $T=722640 426960 1 0 $X=722210 $Y=422405
X266 110 29 28 2 1 2 122 DFFQSRX1 $T=723200 442640 0 0 $X=722770 $Y=442250
X267 126 29 28 2 1 2 139 DFFQSRX1 $T=723200 458320 1 0 $X=722770 $Y=453765
X268 152 29 28 2 1 2 112 DFFQSRX1 $T=758480 395600 0 180 $X=732850 $Y=391045
X269 154 29 28 2 1 2 161 DFFQSRX1 $T=742240 348560 1 0 $X=741810 $Y=344005
X270 155 29 28 2 1 2 169 DFFQSRX1 $T=742240 434800 1 0 $X=741810 $Y=430245
X271 157 29 28 2 1 2 163 DFFQSRX1 $T=742240 442640 1 0 $X=741810 $Y=438085
X272 192 29 28 2 1 2 162 DFFQSRX1 $T=779760 356400 0 180 $X=754130 $Y=351845
X273 188 29 28 2 1 2 166 DFFQSRX1 $T=780880 379920 0 180 $X=755250 $Y=375365
X274 191 29 28 2 1 2 168 DFFQSRX1 $T=781440 379920 1 180 $X=755810 $Y=379530
X275 194 29 28 2 1 2 173 DFFQSRX1 $T=783680 395600 1 180 $X=758050 $Y=395210
X276 185 29 28 2 1 2 178 DFFQSRX1 $T=787040 419120 1 180 $X=761410 $Y=418730
X277 203 29 28 2 1 2 179 DFFQSRX1 $T=792640 411280 1 180 $X=767010 $Y=410890
X278 208 29 28 2 1 2 214 DFFQSRX1 $T=772480 387760 1 0 $X=772050 $Y=383205
X279 220 29 2 28 1 2 222 DFFQSRX1 $T=772480 403440 0 0 $X=772050 $Y=403050
X280 206 29 28 2 1 2 196 DFFQSRX1 $T=797680 426960 1 180 $X=772050 $Y=426570
X281 210 29 28 2 1 2 198 DFFQSRX1 $T=797680 450480 0 180 $X=772050 $Y=445925
X282 35 29 28 2 1 2 22 DFFQSRX1 $T=797680 458320 0 180 $X=772050 $Y=453765
X484 43 42 2 1 41 XOR2X1 $T=629120 442640 1 180 $X=622530 $Y=442250
X485 59 54 2 1 61 XOR2X1 $T=651520 442640 1 0 $X=651090 $Y=438085
X486 56 12 2 1 11 XOR2X1 $T=657680 450480 1 180 $X=651090 $Y=450090
X487 65 60 2 1 67 XOR2X1 $T=663840 426960 0 0 $X=663410 $Y=426570
X488 71 62 2 1 73 XOR2X1 $T=673920 426960 0 0 $X=673490 $Y=426570
X489 82 63 2 1 75 XOR2X1 $T=685120 450480 0 180 $X=678530 $Y=445925
X490 81 79 2 1 84 XOR2X1 $T=684000 426960 1 0 $X=683570 $Y=422405
X491 95 86 2 1 97 XOR2X1 $T=700800 426960 1 0 $X=700370 $Y=422405
X492 96 87 2 1 100 XOR2X1 $T=705840 434800 0 0 $X=705410 $Y=434410
X493 102 106 2 1 101 XOR2X1 $T=731600 419120 0 180 $X=725010 $Y=414565
X494 117 116 2 1 105 XOR2X1 $T=736080 387760 0 180 $X=729490 $Y=383205
X495 123 120 2 1 107 XOR2X1 $T=737760 379920 1 180 $X=731170 $Y=379530
X496 119 121 2 1 109 XOR2X1 $T=737760 419120 1 180 $X=731170 $Y=418730
X497 125 122 2 1 110 XOR2X1 $T=738320 442640 0 180 $X=731730 $Y=438085
X498 137 139 2 1 126 XOR2X1 $T=743920 450480 1 180 $X=737330 $Y=450090
X499 128 135 2 1 115 XOR2X1 $T=745040 364240 0 180 $X=738450 $Y=359685
X500 170 161 2 1 153 XOR2X1 $T=757360 364240 0 180 $X=750770 $Y=359685
X501 160 169 2 1 155 XOR2X1 $T=757920 426960 0 180 $X=751330 $Y=422405
X502 158 18 2 1 17 XOR2X1 $T=758480 458320 0 180 $X=751890 $Y=453765
X503 177 173 2 1 182 XOR2X1 $T=760160 403440 0 0 $X=759730 $Y=403050
X504 176 162 2 1 192 XOR2X1 $T=764080 356400 0 0 $X=763650 $Y=356010
X505 181 178 2 1 183 XOR2X1 $T=765200 419120 1 0 $X=764770 $Y=414565
X506 195 179 2 1 203 XOR2X1 $T=776400 403440 1 0 $X=775970 $Y=398885
X507 204 196 2 1 206 XOR2X1 $T=782000 434800 0 0 $X=781570 $Y=434410
X508 205 198 2 1 210 XOR2X1 $T=787600 442640 1 0 $X=787170 $Y=438085
X509 193 214 2 1 208 XOR2X1 $T=796560 387760 1 180 $X=789970 $Y=387370
X510 229 222 2 1 220 XOR2X1 $T=802160 395600 1 180 $X=795570 $Y=395210
X511 43 42 1 2 3 AND2X1 $T=627440 450480 0 180 $X=623650 $Y=445925
X512 3 4 1 2 5 AND2X1 $T=624080 458320 1 0 $X=623650 $Y=453765
X513 51 46 1 2 43 AND2X1 $T=641440 442640 1 180 $X=637650 $Y=442250
X514 9 53 1 2 56 AND2X1 $T=645360 450480 0 0 $X=644930 $Y=450090
X515 56 12 1 2 59 AND2X1 $T=659360 450480 0 180 $X=655570 $Y=445925
X516 71 62 1 2 65 AND2X1 $T=673360 426960 1 180 $X=669570 $Y=426570
X517 13 73 1 2 74 AND2X1 $T=675600 434800 1 0 $X=675170 $Y=430245
X518 13 75 1 2 76 AND2X1 $T=682880 450480 1 180 $X=679090 $Y=450090
X519 81 77 1 2 71 AND2X1 $T=683440 434800 0 180 $X=679650 $Y=430245
X520 81 79 1 2 82 AND2X1 $T=684560 434800 0 0 $X=684130 $Y=434410
X521 87 86 1 2 85 AND2X1 $T=693520 426960 1 180 $X=689730 $Y=426570
X522 14 15 1 2 91 AND2X1 $T=694640 450480 1 0 $X=694210 $Y=445925
X523 13 94 1 2 16 AND2X1 $T=699680 458320 1 0 $X=699250 $Y=453765
X524 91 89 1 2 96 AND2X1 $T=701920 450480 1 0 $X=701490 $Y=445925
X525 96 87 1 2 95 AND2X1 $T=710320 426960 0 180 $X=706530 $Y=422405
X526 118 115 1 2 113 AND2X1 $T=736640 364240 0 180 $X=732850 $Y=359685
X527 118 107 1 2 114 AND2X1 $T=736640 372080 0 180 $X=732850 $Y=367525
X528 102 106 1 2 119 AND2X1 $T=733280 411280 0 0 $X=732850 $Y=410890
X529 108 111 1 2 102 AND2X1 $T=737200 403440 1 180 $X=733410 $Y=403050
X530 117 116 1 2 123 AND2X1 $T=741120 387760 0 180 $X=737330 $Y=383205
X531 125 122 1 2 137 AND2X1 $T=738880 442640 1 0 $X=738450 $Y=438085
X532 138 140 1 2 124 AND2X1 $T=745600 372080 0 180 $X=741810 $Y=367525
X533 146 112 1 2 108 AND2X1 $T=747280 403440 1 180 $X=743490 $Y=403050
X534 106 121 1 2 148 AND2X1 $T=743920 419120 1 0 $X=743490 $Y=414565
X535 118 151 1 2 152 AND2X1 $T=748400 403440 1 0 $X=747970 $Y=398885
X536 118 153 1 2 154 AND2X1 $T=754560 356400 0 180 $X=750770 $Y=351845
X537 165 163 1 2 158 AND2X1 $T=761840 450480 0 180 $X=758050 $Y=445925
X538 176 162 1 2 170 AND2X1 $T=762960 356400 1 180 $X=759170 $Y=356010
X539 158 18 1 2 19 AND2X1 $T=759600 458320 1 0 $X=759170 $Y=453765
X540 160 169 1 2 181 AND2X1 $T=761280 426960 1 0 $X=760850 $Y=422405
X541 160 174 1 2 177 AND2X1 $T=761840 419120 1 0 $X=761410 $Y=414565
X542 168 166 1 2 176 AND2X1 $T=762960 372080 1 0 $X=762530 $Y=367525
X543 118 183 1 2 185 AND2X1 $T=764080 411280 0 0 $X=763650 $Y=410890
X544 118 182 1 2 194 AND2X1 $T=768000 403440 0 0 $X=767570 $Y=403050
X545 177 173 1 2 195 AND2X1 $T=769120 403440 1 0 $X=768690 $Y=398885
X546 204 196 1 2 205 AND2X1 $T=782560 442640 1 0 $X=782130 $Y=438085
X547 23 202 1 2 204 AND2X1 $T=783120 450480 0 0 $X=782690 $Y=450090
X548 28 209 1 2 215 AND2X1 $T=798240 364240 0 180 $X=794450 $Y=359685
X549 233 234 1 2 211 AND2X1 $T=798800 332880 1 0 $X=798370 $Y=328325
X550 28 241 1 2 231 AND2X1 $T=805520 372080 0 180 $X=801730 $Y=367525
X551 251 246 1 2 243 AND2X1 $T=807200 317200 1 180 $X=803410 $Y=316810
X552 259 254 1 2 252 AND2X1 $T=810560 348560 0 180 $X=806770 $Y=344005
X553 28 264 1 2 248 AND2X1 $T=810000 372080 0 0 $X=809570 $Y=371690
X554 222 269 1 2 274 AND2X1 $T=812240 387760 1 0 $X=811810 $Y=383205
X555 283 289 1 2 287 AND2X1 $T=819520 387760 1 0 $X=819090 $Y=383205
X556 265 261 1 2 233 AND2X1 $T=825120 340720 1 180 $X=821330 $Y=340330
X590 42 44 1 2 45 OR2X1 $T=629120 442640 0 0 $X=628690 $Y=442250
X591 4 45 1 2 7 OR2X1 $T=629680 458320 1 0 $X=629250 $Y=453765
X592 46 50 1 2 44 OR2X1 $T=636400 450480 0 180 $X=632610 $Y=445925
X593 54 57 1 2 50 OR2X1 $T=650960 442640 1 180 $X=647170 $Y=442250
X594 12 64 1 2 57 OR2X1 $T=659360 450480 1 0 $X=658930 $Y=445925
X595 60 66 1 2 64 OR2X1 $T=667200 442640 0 180 $X=663410 $Y=438085
X596 86 88 1 2 83 OR2X1 $T=695760 434800 1 180 $X=691970 $Y=434410
X597 122 129 1 2 133 OR2X1 $T=737760 434800 1 0 $X=737330 $Y=430245
X598 111 131 1 2 132 OR2X1 $T=738880 403440 0 0 $X=738450 $Y=403050
X599 106 132 1 2 136 OR2X1 $T=738880 411280 0 0 $X=738450 $Y=410890
X600 121 136 1 2 129 OR2X1 $T=743360 419120 1 180 $X=739570 $Y=418730
X601 139 133 1 2 145 OR2X1 $T=743360 434800 0 0 $X=742930 $Y=434410
X602 150 130 1 2 149 OR2X1 $T=750640 372080 1 180 $X=746850 $Y=371690
X603 169 145 1 2 175 OR2X1 $T=762400 434800 1 180 $X=758610 $Y=434410
X604 163 175 1 2 180 OR2X1 $T=766880 450480 0 180 $X=763090 $Y=445925
X605 18 180 1 2 20 OR2X1 $T=766880 458320 0 180 $X=763090 $Y=453765
X606 168 184 1 2 118 OR2X1 $T=768000 387760 1 180 $X=764210 $Y=387370
X607 179 186 1 2 184 OR2X1 $T=769120 411280 0 180 $X=765330 $Y=406725
X608 198 24 1 2 200 OR2X1 $T=779200 434800 1 180 $X=775410 $Y=434410
X609 26 243 1 2 247 OR2X1 $T=802160 325040 1 0 $X=801730 $Y=320485
X610 261 257 1 2 218 OR2X1 $T=811120 340720 1 180 $X=807330 $Y=340330
X611 272 267 1 2 255 OR2X1 $T=815040 356400 0 180 $X=811250 $Y=351845
X612 253 269 1 2 277 OR2X1 $T=815040 364240 0 0 $X=814610 $Y=363850
X613 280 261 1 2 272 OR2X1 $T=818960 325040 0 180 $X=815170 $Y=320485
X614 261 267 1 2 295 OR2X1 $T=821200 356400 1 0 $X=820770 $Y=351845
X615 282 293 1 2 299 OR2X1 $T=823440 395600 1 0 $X=823010 $Y=391045
X616 282 296 1 2 292 OR2X1 $T=826800 403440 1 180 $X=823010 $Y=403050
X617 276 299 1 2 291 OR2X1 $T=824560 395600 0 0 $X=824130 $Y=395210
X618 6 46 42 1 2 47 NAND3X1 $T=630240 450480 0 0 $X=629810 $Y=450090
X619 52 54 12 1 2 58 NAND3X1 $T=652080 450480 1 0 $X=651650 $Y=445925
X620 70 60 62 1 2 68 NAND3X1 $T=672800 442640 0 180 $X=668450 $Y=438085
X621 72 62 63 1 2 66 NAND3X1 $T=677840 442640 0 180 $X=673490 $Y=438085
X622 85 15 89 1 2 80 NAND3X1 $T=691840 442640 1 0 $X=691410 $Y=438085
X623 92 93 15 1 2 88 NAND3X1 $T=700800 434800 1 180 $X=696450 $Y=434410
X624 142 112 120 1 2 131 NAND3X1 $T=745600 387760 0 180 $X=741250 $Y=383205
X625 143 120 116 1 2 141 NAND3X1 $T=746720 379920 1 180 $X=742370 $Y=379530
X626 148 112 111 1 2 147 NAND3X1 $T=748400 411280 0 180 $X=744050 $Y=406725
X627 164 161 135 1 2 150 NAND3X1 $T=756240 372080 0 180 $X=751890 $Y=367525
X628 176 162 161 1 2 138 NAND3X1 $T=760720 364240 1 180 $X=756370 $Y=363850
X629 171 179 173 1 2 167 NAND3X1 $T=760160 411280 1 0 $X=759730 $Y=406725
X630 21 163 18 1 2 187 NAND3X1 $T=769680 450480 1 180 $X=765330 $Y=450090
X631 199 173 178 1 2 186 NAND3X1 $T=775840 419120 0 180 $X=771490 $Y=414565
X632 201 198 196 1 2 197 NAND3X1 $T=776400 442640 0 0 $X=775970 $Y=442250
X633 213 223 228 1 2 225 NAND3X1 $T=795440 348560 1 0 $X=795010 $Y=344005
X634 255 252 238 1 2 236 NAND3X1 $T=810000 348560 1 180 $X=805650 $Y=348170
X635 258 253 242 1 2 251 NAND3X1 $T=810560 325040 1 180 $X=806210 $Y=324650
X636 233 257 249 1 2 254 NAND3X1 $T=811680 332880 1 180 $X=807330 $Y=332490
X637 263 261 268 1 2 224 NAND3X1 $T=810560 317200 1 0 $X=810130 $Y=312645
X638 263 261 260 1 2 259 NAND3X1 $T=814480 325040 0 180 $X=810130 $Y=320485
X639 272 253 265 1 2 228 NAND3X1 $T=816160 348560 0 180 $X=811810 $Y=344005
X640 267 275 277 1 2 278 NAND3X1 $T=815040 356400 0 0 $X=814610 $Y=356010
X641 262 265 286 1 2 275 NAND3X1 $T=816160 356400 1 0 $X=815730 $Y=351845
X642 287 279 266 1 2 270 NAND3X1 $T=820640 403440 1 180 $X=816290 $Y=403050
X643 263 242 280 1 2 290 NAND3X1 $T=818960 325040 1 0 $X=818530 $Y=320485
X644 287 288 297 1 2 296 NAND3X1 $T=821200 403440 1 0 $X=820770 $Y=398885
X645 285 271 265 1 2 298 NAND3X1 $T=822320 332880 1 0 $X=821890 $Y=328325
X646 247 290 298 1 2 300 NAND3X1 $T=823440 325040 1 0 $X=823010 $Y=320485
X647 301 295 302 1 2 303 NAND3X1 $T=826240 348560 0 0 $X=825810 $Y=348170
X648 49 43 1 2 48 NOR2X1 $T=635280 442640 1 180 $X=632050 $Y=442250
X649 46 51 1 2 49 NOR2X1 $T=640880 442640 0 180 $X=637650 $Y=438085
X650 8 47 1 2 52 NOR2X1 $T=641440 450480 1 180 $X=638210 $Y=450090
X651 47 55 1 2 9 NOR2X1 $T=643120 450480 1 0 $X=642690 $Y=445925
X652 58 55 1 2 10 NOR2X1 $T=651520 450480 1 180 $X=648290 $Y=450090
X653 69 68 1 2 51 NOR2X1 $T=672240 450480 0 180 $X=669010 $Y=445925
X654 78 80 1 2 70 NOR2X1 $T=680080 442640 1 0 $X=679650 $Y=438085
X655 80 69 1 2 81 NOR2X1 $T=686240 442640 0 0 $X=685810 $Y=442250
X656 79 83 1 2 72 NOR2X1 $T=686800 434800 1 0 $X=686370 $Y=430245
X657 15 14 1 2 90 NOR2X1 $T=695200 458320 1 0 $X=694770 $Y=453765
X658 90 91 1 2 94 NOR2X1 $T=699680 450480 0 0 $X=699250 $Y=450090
X659 89 91 1 2 98 NOR2X1 $T=705280 450480 0 0 $X=704850 $Y=450090
X660 98 96 1 2 99 NOR2X1 $T=708080 450480 1 0 $X=707650 $Y=445925
X661 104 102 1 2 103 NOR2X1 $T=730480 403440 1 180 $X=727250 $Y=403050
X662 111 108 1 2 104 NOR2X1 $T=733840 403440 1 180 $X=730610 $Y=403050
X663 124 128 1 2 127 NOR2X1 $T=736640 356400 0 0 $X=736210 $Y=356010
X664 134 138 1 2 117 NOR2X1 $T=740000 379920 0 0 $X=739570 $Y=379530
X665 112 146 1 2 144 NOR2X1 $T=744480 403440 1 0 $X=744050 $Y=398885
X666 140 138 1 2 128 NOR2X1 $T=747280 364240 1 0 $X=746850 $Y=359685
X667 116 149 1 2 142 NOR2X1 $T=747280 387760 0 0 $X=746850 $Y=387370
X668 138 141 1 2 146 NOR2X1 $T=751760 379920 1 180 $X=748530 $Y=379530
X669 144 108 1 2 151 NOR2X1 $T=748960 403440 0 0 $X=748530 $Y=403050
X670 156 158 1 2 157 NOR2X1 $T=751200 450480 1 0 $X=750770 $Y=445925
X671 147 159 1 2 160 NOR2X1 $T=752320 411280 0 0 $X=751890 $Y=410890
X672 159 167 1 2 165 NOR2X1 $T=754000 419120 1 0 $X=753570 $Y=414565
X673 163 165 1 2 156 NOR2X1 $T=754000 450480 1 0 $X=753570 $Y=445925
X674 172 147 1 2 171 NOR2X1 $T=757920 411280 0 180 $X=754690 $Y=406725
X675 162 166 1 2 164 NOR2X1 $T=758480 372080 1 0 $X=758050 $Y=367525
X676 190 176 1 2 188 NOR2X1 $T=769120 364240 1 180 $X=765890 $Y=363850
X677 168 193 1 2 191 NOR2X1 $T=768000 387760 0 0 $X=767570 $Y=387370
X678 166 168 1 2 190 NOR2X1 $T=771360 372080 0 180 $X=768130 $Y=367525
X679 197 189 1 2 125 NOR2X1 $T=773600 442640 0 180 $X=770370 $Y=438085
X680 187 189 1 2 23 NOR2X1 $T=774720 450480 1 180 $X=771490 $Y=450090
X681 25 187 1 2 201 NOR2X1 $T=779200 450480 1 180 $X=775970 $Y=450090
X682 196 200 1 2 199 NOR2X1 $T=782000 434800 1 180 $X=778770 $Y=434410
X683 207 216 1 2 212 NOR2X1 $T=793760 325040 1 0 $X=793330 $Y=320485
X684 211 217 1 2 213 NOR2X1 $T=793760 332880 1 0 $X=793330 $Y=328325
X685 218 221 1 2 219 NOR2X1 $T=794880 340720 1 0 $X=794450 $Y=336165
X686 27 224 1 2 217 NOR2X1 $T=796000 317200 1 0 $X=795570 $Y=312645
X687 27 216 1 2 227 NOR2X1 $T=797680 317200 0 0 $X=797250 $Y=316810
X688 230 219 1 2 223 NOR2X1 $T=800480 340720 0 180 $X=797250 $Y=336165
X689 226 232 1 2 229 NOR2X1 $T=797680 395600 1 0 $X=797250 $Y=391045
X690 212 227 1 2 221 NOR2X1 $T=798240 325040 0 0 $X=797810 $Y=324650
X691 244 26 1 2 237 NOR2X1 $T=804960 340720 1 180 $X=801730 $Y=340330
X692 237 218 1 2 235 NOR2X1 $T=802160 348560 1 0 $X=801730 $Y=344005
X693 240 245 1 2 230 NOR2X1 $T=802720 340720 1 0 $X=802290 $Y=336165
X694 244 272 1 2 258 NOR2X1 $T=813360 332880 0 0 $X=812930 $Y=332490
X695 253 272 1 2 273 NOR2X1 $T=813360 340720 1 0 $X=812930 $Y=336165
X696 268 261 1 2 256 NOR2X1 $T=814480 317200 1 0 $X=814050 $Y=312645
X697 265 253 1 2 263 NOR2X1 $T=818960 348560 0 180 $X=815730 $Y=344005
X698 242 285 1 2 281 NOR2X1 $T=817840 332880 1 0 $X=817410 $Y=328325
X699 273 281 1 2 245 NOR2X1 $T=817840 340720 1 0 $X=817410 $Y=336165
X700 31 240 1 2 282 NOR2X1 $T=820640 372080 1 180 $X=817410 $Y=371690
X701 253 284 1 2 294 NOR2X1 $T=824560 332880 1 180 $X=821330 $Y=332490
X702 31 253 1 2 276 NOR2X1 $T=826240 372080 1 180 $X=823010 $Y=371690
X703 294 300 1 2 301 NOR2X1 $T=826800 332880 0 0 $X=826370 $Y=332490
X734 8 1 2 53 INVX2 $T=640880 458320 1 0 $X=640450 $Y=453765
X735 51 1 2 55 INVX2 $T=643680 442640 0 0 $X=643250 $Y=442250
X736 78 1 2 77 INVX2 $T=681760 426960 1 180 $X=679650 $Y=426570
X737 14 1 2 69 INVX2 $T=689600 450480 0 180 $X=687490 $Y=445925
X738 89 1 2 92 INVX2 $T=697440 442640 0 0 $X=697010 $Y=442250
X739 87 1 2 93 INVX2 $T=702480 434800 1 180 $X=700370 $Y=434410
X740 134 1 2 143 INVX2 $T=747280 379920 0 180 $X=745170 $Y=375365
X741 130 1 2 140 INVX2 $T=748400 364240 0 0 $X=747970 $Y=363850
X742 146 1 2 159 INVX2 $T=752320 411280 1 0 $X=751890 $Y=406725
X743 172 1 2 174 INVX2 $T=757920 411280 0 0 $X=757490 $Y=410890
X744 165 1 2 189 INVX2 $T=766880 450480 1 0 $X=766450 $Y=445925
X745 118 1 2 193 INVX2 $T=770800 395600 1 0 $X=770370 $Y=391045
X746 25 1 2 202 INVX2 $T=779200 450480 0 0 $X=778770 $Y=450090
X747 26 1 2 207 INVX2 $T=789280 325040 1 0 $X=788850 $Y=320485
X748 214 1 2 232 INVX2 $T=800480 387760 0 0 $X=800050 $Y=387370
X749 27 1 2 242 INVX2 $T=802720 317200 1 0 $X=802290 $Y=312645
X750 218 1 2 262 INVX2 $T=810000 348560 0 0 $X=809570 $Y=348170
X751 31 1 2 28 INVX2 $T=810560 387760 1 0 $X=810130 $Y=383205
X752 253 1 2 257 INVX2 $T=811680 332880 1 0 $X=811250 $Y=328325
X753 244 1 2 249 INVX2 $T=813360 332880 1 180 $X=811250 $Y=332490
X754 261 1 2 269 INVX2 $T=813920 372080 0 0 $X=813490 $Y=371690
X755 276 1 2 279 INVX2 $T=817280 395600 0 0 $X=816850 $Y=395210
X756 281 1 2 284 INVX2 $T=818400 332880 0 0 $X=817970 $Y=332490
X757 240 1 2 265 INVX2 $T=818960 348560 1 0 $X=818530 $Y=344005
X758 256 1 2 285 INVX2 $T=819520 317200 1 0 $X=819090 $Y=312645
X759 268 1 2 280 INVX2 $T=825120 317200 1 180 $X=823010 $Y=316810
X782 79 63 1 2 78 NAND2X1 $T=682880 434800 1 180 $X=679650 $Y=434410
X783 130 135 1 2 134 NAND2X1 $T=739440 372080 1 0 $X=739010 $Y=367525
X784 169 178 1 2 172 NAND2X1 $T=759040 419120 0 0 $X=758610 $Y=418730
X785 235 240 1 2 238 NAND2X1 $T=801600 348560 0 0 $X=801170 $Y=348170
X786 242 26 1 2 239 NAND2X1 $T=804960 325040 1 180 $X=801730 $Y=324650
X787 239 249 1 2 234 NAND2X1 $T=803280 332880 1 0 $X=802850 $Y=328325
X788 240 249 1 2 216 NAND2X1 $T=805520 340720 1 0 $X=805090 $Y=336165
X789 227 256 1 2 246 NAND2X1 $T=807200 317200 0 0 $X=806770 $Y=316810
X790 30 31 1 2 266 NAND2X1 $T=811680 411280 1 0 $X=811250 $Y=406725
X791 242 268 1 2 260 NAND2X1 $T=812800 317200 0 0 $X=812370 $Y=316810
X792 257 242 1 2 271 NAND2X1 $T=813360 332880 1 0 $X=812930 $Y=328325
X793 274 28 1 2 283 NAND2X1 $T=817840 387760 0 0 $X=817410 $Y=387370
X794 276 261 1 2 288 NAND2X1 $T=819520 395600 1 0 $X=819090 $Y=391045
X795 263 286 1 2 267 NAND2X1 $T=820080 348560 0 0 $X=819650 $Y=348170
X796 282 261 1 2 289 NAND2X1 $T=820080 379920 0 0 $X=819650 $Y=379530
X797 233 244 1 2 302 NAND2X1 $T=826800 348560 1 0 $X=826370 $Y=344005
X798 33 31 1 2 297 NAND2X1 $T=831280 403440 0 180 $X=828050 $Y=398885
X826 29 209 2 225 1 DFFQX1 $T=803280 356400 0 180 $X=790530 $Y=351845
X827 29 240 2 231 1 DFFQX1 $T=797680 372080 0 0 $X=797250 $Y=371690
X828 29 253 2 215 1 DFFQX1 $T=800480 364240 1 0 $X=800050 $Y=359685
X829 29 264 2 236 1 DFFQX1 $T=800480 364240 0 0 $X=800050 $Y=363850
X830 29 261 2 248 1 DFFQX1 $T=803280 379920 0 0 $X=802850 $Y=379530
X831 29 226 2 250 1 DFFQX1 $T=815600 395600 1 180 $X=802850 $Y=395210
X832 29 30 2 270 1 DFFQX1 $T=816160 411280 1 180 $X=803410 $Y=410890
X833 29 32 2 291 1 DFFQX1 $T=820080 411280 1 0 $X=819650 $Y=406725
X834 29 33 2 292 1 DFFQX1 $T=820080 419120 1 0 $X=819650 $Y=414565
X835 29 286 2 278 1 DFFQX1 $T=832960 356400 1 180 $X=820210 $Y=356010
X836 29 241 2 303 1 DFFQX1 $T=832960 364240 1 180 $X=820210 $Y=363850
X853 214 31 226 1 2 250 MUX2X1 $T=811120 387760 1 180 $X=805090 $Y=387370
X854 32 28 274 1 2 293 MUX2X1 $T=828480 387760 0 180 $X=822450 $Y=383205
.ENDS
***************************************
.SUBCKT ICV_43
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_45
** N=5 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_46
** N=7 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT ICV_47
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39
** N=4 EP=0 IP=16 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_41
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_42
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_49 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 27 28 29 30 31 32 35
** N=172 EP=32 IP=1889 FDC=1504
M0 1 40 2 1 N L=1.8e-07 W=2.2e-07 $X=625400 $Y=482600 $D=0
M1 3 40 2 3 P L=1.8e-07 W=4.4e-07 $X=625400 $Y=484555 $D=16
X2 3 1 35 1 pad_out $T=1726400 503200 0 90 $X=1492300 $Y=502300
X90 41 28 2 3 1 3 4 DFFQSRX1 $T=611760 466160 0 0 $X=611330 $Y=465770
X91 27 28 29 3 1 3 40 DFFQSRX1 $T=612320 489680 0 0 $X=611890 $Y=489290
X92 42 28 2 3 1 3 43 DFFQSRX1 $T=612880 481840 1 0 $X=612450 $Y=477285
X93 53 28 2 3 1 3 46 DFFQSRX1 $T=664960 481840 1 180 $X=639330 $Y=481450
X94 30 28 2 3 1 3 12 DFFQSRX1 $T=640880 458320 0 0 $X=640450 $Y=457930
X95 54 28 2 3 1 3 45 DFFQSRX1 $T=666080 474000 0 180 $X=640450 $Y=469445
X96 55 28 2 3 1 3 48 DFFQSRX1 $T=667200 489680 0 180 $X=641570 $Y=485125
X97 56 28 2 3 1 3 49 DFFQSRX1 $T=667200 505360 0 180 $X=641570 $Y=500805
X98 66 28 2 3 1 3 69 DFFQSRX1 $T=657680 497520 0 0 $X=657250 $Y=497130
X99 63 28 2 3 1 3 62 DFFQSRX1 $T=666080 474000 1 0 $X=665650 $Y=469445
X100 73 28 2 3 1 3 58 DFFQSRX1 $T=693520 466160 1 180 $X=667890 $Y=465770
X101 31 28 2 3 1 3 15 DFFQSRX1 $T=689040 458320 0 0 $X=688610 $Y=457930
X102 79 28 2 3 1 3 76 DFFQSRX1 $T=689040 505360 0 0 $X=688610 $Y=504970
X103 93 28 2 3 1 3 85 DFFQSRX1 $T=724320 466160 1 180 $X=698690 $Y=465770
X104 92 28 2 3 1 3 84 DFFQSRX1 $T=724320 474000 1 180 $X=698690 $Y=473610
X105 94 28 2 3 1 3 86 DFFQSRX1 $T=725440 497520 1 180 $X=699810 $Y=497130
X106 97 28 2 3 1 3 88 DFFQSRX1 $T=739440 481840 0 180 $X=713810 $Y=477285
X107 96 28 2 3 1 3 98 DFFQSRX1 $T=715920 489680 1 0 $X=715490 $Y=485125
X108 32 28 29 3 1 3 18 DFFQSRX1 $T=743360 458320 0 0 $X=742930 $Y=457930
X109 102 28 29 3 1 3 105 DFFQSRX1 $T=745040 474000 0 0 $X=744610 $Y=473610
X110 104 28 29 3 1 3 106 DFFQSRX1 $T=746160 489680 1 0 $X=745730 $Y=485125
X111 119 28 29 3 1 3 114 DFFQSRX1 $T=797680 474000 1 180 $X=772050 $Y=473610
X112 120 28 29 3 1 3 25 DFFQSRX1 $T=772480 489680 0 0 $X=772050 $Y=489290
X199 5 4 3 1 41 XOR2X1 $T=628000 458320 1 180 $X=621410 $Y=457930
X200 6 43 3 1 42 XOR2X1 $T=629120 474000 0 180 $X=622530 $Y=469445
X201 51 46 3 1 53 XOR2X1 $T=648160 474000 0 0 $X=647730 $Y=473610
X202 10 45 3 1 54 XOR2X1 $T=650960 466160 1 0 $X=650530 $Y=461605
X203 11 48 3 1 55 XOR2X1 $T=650960 497520 1 0 $X=650530 $Y=492965
X204 52 49 3 1 56 XOR2X1 $T=651520 513200 1 0 $X=651090 $Y=508645
X205 64 62 3 1 59 XOR2X1 $T=680080 481840 1 180 $X=673490 $Y=481450
X206 67 58 3 1 73 XOR2X1 $T=679520 466160 1 0 $X=679090 $Y=461605
X207 75 69 3 1 68 XOR2X1 $T=690160 497520 0 180 $X=683570 $Y=492965
X208 89 86 3 1 91 XOR2X1 $T=704720 497520 1 0 $X=704290 $Y=492965
X209 87 85 3 1 93 XOR2X1 $T=708080 481840 0 0 $X=707650 $Y=481450
X210 95 98 3 1 96 XOR2X1 $T=731040 497520 0 180 $X=724450 $Y=492965
X211 107 105 3 1 102 XOR2X1 $T=762400 466160 1 180 $X=755810 $Y=465770
X212 16 106 3 1 104 XOR2X1 $T=762960 481840 0 180 $X=756370 $Y=477285
X213 108 101 3 1 103 XOR2X1 $T=764080 497520 0 180 $X=757490 $Y=492965
X214 111 112 3 1 117 XOR2X1 $T=769120 505360 1 0 $X=768690 $Y=500805
X215 23 114 3 1 119 XOR2X1 $T=782560 466160 0 0 $X=782130 $Y=465770
X216 118 21 3 1 24 XOR2X1 $T=788160 466160 1 0 $X=787730 $Y=461605
X217 4 43 1 3 7 AND2X1 $T=633600 458320 1 180 $X=629810 $Y=457930
X218 10 45 1 3 51 AND2X1 $T=645920 466160 1 0 $X=645490 $Y=461605
X219 11 48 1 3 52 AND2X1 $T=654880 497520 1 180 $X=651090 $Y=497130
X220 13 59 1 3 63 AND2X1 $T=680640 481840 0 180 $X=676850 $Y=477285
X221 13 68 1 3 66 AND2X1 $T=682880 497520 0 180 $X=679090 $Y=492965
X222 67 58 1 3 64 AND2X1 $T=683440 481840 1 180 $X=679650 $Y=481450
X223 77 78 1 3 80 AND2X1 $T=694640 497520 1 0 $X=694210 $Y=492965
X224 88 84 1 3 87 AND2X1 $T=703600 481840 0 180 $X=699810 $Y=477285
X225 87 85 1 3 89 AND2X1 $T=709200 489680 0 180 $X=705410 $Y=485125
X226 13 91 1 3 94 AND2X1 $T=712000 497520 1 0 $X=711570 $Y=492965
X227 16 106 1 3 107 AND2X1 $T=762960 481840 1 0 $X=762530 $Y=477285
X228 106 105 1 3 19 AND2X1 $T=765760 466160 1 0 $X=765330 $Y=461605
X229 23 114 1 3 118 AND2X1 $T=782560 466160 1 0 $X=782130 $Y=461605
X230 43 8 1 3 44 OR2X1 $T=630240 474000 1 0 $X=629810 $Y=469445
X231 45 44 1 3 47 OR2X1 $T=637520 474000 1 0 $X=637090 $Y=469445
X232 46 47 1 3 50 OR2X1 $T=643680 474000 0 0 $X=643250 $Y=473610
X233 88 61 1 3 13 OR2X1 $T=703040 497520 0 180 $X=699250 $Y=492965
X234 105 17 1 3 109 OR2X1 $T=763520 466160 0 0 $X=763090 $Y=465770
X235 106 109 1 3 113 OR2X1 $T=769120 466160 0 0 $X=768690 $Y=465770
X236 112 110 1 3 116 OR2X1 $T=771920 497520 1 0 $X=771490 $Y=492965
X237 21 115 1 3 20 OR2X1 $T=777520 458320 1 180 $X=773730 $Y=457930
X238 114 113 1 3 115 OR2X1 $T=777520 466160 0 180 $X=773730 $Y=461605
X239 57 60 62 1 3 61 NAND3X1 $T=673920 497520 1 0 $X=673490 $Y=492965
X240 72 62 58 1 3 70 NAND3X1 $T=685680 481840 0 180 $X=681330 $Y=477285
X241 82 83 86 1 3 81 NAND3X1 $T=696320 481840 0 0 $X=695890 $Y=481450
X242 87 85 86 1 3 77 NAND3X1 $T=704720 489680 0 180 $X=700370 $Y=485125
X243 48 49 1 3 57 NOR2X1 $T=657120 497520 1 0 $X=656690 $Y=492965
X244 58 65 1 3 60 NOR2X1 $T=677840 489680 1 0 $X=677410 $Y=485125
X245 77 70 1 3 14 NOR2X1 $T=691280 481840 0 180 $X=688050 $Y=477285
X246 74 77 1 3 67 NOR2X1 $T=688480 481840 0 0 $X=688050 $Y=481450
X247 80 75 1 3 79 NOR2X1 $T=692960 497520 0 180 $X=689730 $Y=492965
X248 76 81 1 3 71 NOR2X1 $T=692960 489680 1 0 $X=692530 $Y=485125
X249 78 77 1 3 75 NOR2X1 $T=695200 489680 0 0 $X=694770 $Y=489290
X250 84 50 1 3 82 NOR2X1 $T=699680 481840 0 180 $X=696450 $Y=477285
X251 84 88 1 3 90 NOR2X1 $T=705840 481840 1 0 $X=705410 $Y=477285
X252 90 87 1 3 92 NOR2X1 $T=709760 481840 1 0 $X=709330 $Y=477285
X253 88 95 1 3 97 NOR2X1 $T=724880 481840 0 0 $X=724450 $Y=481450
X258 74 1 3 72 INVX2 $T=686240 481840 0 0 $X=685810 $Y=481450
X259 76 1 3 78 INVX2 $T=691840 489680 1 180 $X=689730 $Y=489290
X260 85 1 3 83 INVX2 $T=704720 481840 1 180 $X=702610 $Y=481450
X261 13 1 3 95 INVX2 $T=717600 497520 1 0 $X=717170 $Y=492965
X262 98 1 3 99 INVX2 $T=736640 497520 1 0 $X=736210 $Y=492965
X263 101 1 3 100 INVX2 $T=750080 489680 1 180 $X=747970 $Y=489290
X264 110 1 3 111 INVX2 $T=772480 497520 1 180 $X=770370 $Y=497130
X265 45 46 1 3 9 NAND2X1 $T=641440 466160 1 0 $X=641010 $Y=461605
X266 71 69 1 3 65 NAND2X1 $T=682880 489680 1 0 $X=682450 $Y=485125
X267 76 69 1 3 74 NAND2X1 $T=690720 489680 0 180 $X=687490 $Y=485125
X268 108 101 1 3 110 NAND2X1 $T=769120 497520 0 180 $X=765890 $Y=492965
X269 114 21 1 3 22 NAND2X1 $T=777520 466160 1 0 $X=777090 $Y=461605
X277 99 101 3 100 1 DFFQX1 $T=742800 497520 0 0 $X=742370 $Y=497130
X278 99 108 3 103 1 DFFQX1 $T=754560 505360 1 0 $X=754130 $Y=500805
X279 99 112 3 117 1 DFFQX1 $T=776400 505360 1 0 $X=775970 $Y=500805
X280 99 120 3 116 1 DFFQX1 $T=778080 497520 0 0 $X=777650 $Y=497130
.ENDS
***************************************
.SUBCKT ICV_19
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=7 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=19 EP=0 IP=22 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=35 EP=0 IP=38 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 5 7 8
** N=63 EP=5 IP=1047 FDC=192
X0 2 1 7 1 pad_out $T=1726400 683200 0 90 $X=1492300 $Y=682300
X1 2 5 8 1 pad_out $T=1726400 773200 0 90 $X=1492300 $Y=772300
.ENDS
***************************************
.SUBCKT ICV_26 1 2 6 7 8
** N=63 EP=5 IP=1047 FDC=192
X0 2 1 7 1 pad_out $T=1726400 863200 0 90 $X=1492300 $Y=862300
X1 2 6 8 1 pad_out $T=1726400 953200 0 90 $X=1492300 $Y=952300
.ENDS
***************************************
.SUBCKT ICV_25 1 2 6 7
** N=73 EP=4 IP=1506 FDC=192
X0 2 1 6 1 pad_out $T=1726400 1133200 0 90 $X=1492300 $Y=1132300
X1 2 1 7 1 pad_out $T=1726400 1223200 0 90 $X=1492300 $Y=1222300
.ENDS
***************************************
.SUBCKT ICV_2 VSS VDD
** N=46 EP=2 IP=1 FDC=1
D0 VSS VDD ndio_m AREA=9e-10 PJ=0.00012 $X=10780 $Y=193610 $D=30
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3
** N=5 EP=3 IP=6 FDC=96
X0 2 1 3 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4
** N=6 EP=4 IP=6 FDC=96
X0 2 3 4 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3
** N=5 EP=3 IP=6 FDC=96
X0 2 1 3 1 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT soc_top VSS VDD clk h0_4 h0_0 h1_5 h1_1 m0_5 m0_1 m1_6 m1_2 s0_6 s0_2 s1_3 btn_light h0_3 colon h1_4 h1_0 m0_4
+ m0_0 m1_5 m1_1 s0_5 s0_1 s1_6 s1_2 s1_5 btn_mode btn_dec h0_5 h0_1 h1_6 h1_2 m0_6 m0_2 reset m1_3 s1_0 s0_3
+ s1_4 btn_set btn_inc h0_2 h1_3 m1_0 m0_3 s0_0 s1_1 s0_4 h0_6 light m1_4
** N=94 EP=53 IP=231 FDC=9126
X1 VSS VDD 22 clk h0_4 ICV_69 $T=0 0 0 0 $X=0 $Y=232300
X2 VSS VDD 4 h0_0 ICV_8 $T=0 503200 0 270 $X=0 $Y=412300
X4 VSS VDD ICV_1 $T=0 593200 0 270 $X=0 $Y=502300
X5 VSS VDD h1_5 ICV_6 $T=0 683200 0 270 $X=0 $Y=592300
X6 VSS VDD h1_1 m0_5 ICV_67 $T=0 0 0 0 $X=0 $Y=680200
X7 VSS VDD m0_1 m1_6 ICV_66 $T=0 0 0 0 $X=0 $Y=862300
X8 VSS VDD m1_2 ICV_4 $T=0 1133200 0 270 $X=0 $Y=1042300
X9 VSS VDD s0_6 s0_2 ICV_65 $T=0 0 0 0 $X=0 $Y=1130200
X10 VSS VDD s1_3 ICV_64 $T=0 0 0 0 $X=0 $Y=1312300
X11 VSS VDD 3 4 5 btn_light h0_3 colon h1_4 h1_0 m0_4 m0_0 m1_5 m1_1 s0_5 s0_1 s1_6 s1_2 s1_5 ICV_9 $T=0 0 0 0 $X=232300 $Y=1312300
X12 VSS VDD 6 7 8 9 btn_mode btn_dec reset h0_5 h0_1 h1_6 h1_2 m0_6 m0_2 m1_3 s1_0 s0_3 s1_4 ICV_63 $T=0 0 0 0 $X=232600 $Y=0
X13 VSS VDD 10 11 12 13 14 15 16 30 23 24 32 33 17 25 26 18 27 28
+ 19 20 37 35 36 7 6 34 22 4 8 9 5 31 21 btn_set btn_inc
+ ICV_59 $T=0 0 0 0 $X=234100 $Y=232300
X14 VSS 31 VDD 11 10 12 13 14 15 16 30 24 32 33 17 27 28 18 19 35
+ 20 36 37 21 29 3 22 34 23 25 26 h0_2
+ ICV_49 $T=0 0 0 0 $X=234100 $Y=457930
X15 VSS VDD 5 h1_3 m1_0 ICV_27 $T=0 0 0 0 $X=234100 $Y=665400
X16 VSS VDD 9 m0_3 s0_0 ICV_26 $T=0 0 0 0 $X=234100 $Y=862300
X17 VSS VDD s1_1 s0_4 ICV_25 $T=0 0 0 0 $X=234100 $Y=1073125
X18 VSS VDD ICV_2 $T=413200 1636400 0 180 $X=322300 $Y=1402300
X19 VSS VDD h0_6 ICV_7 $T=1726400 413200 0 90 $X=1492300 $Y=412300
X20 VSS VDD 29 light ICV_5 $T=1726400 593200 0 90 $X=1492300 $Y=592300
X21 VSS VDD m1_4 ICV_3 $T=1726400 1043200 0 90 $X=1492300 $Y=1042300
.ENDS
***************************************

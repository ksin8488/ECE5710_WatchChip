* SPICE NETLIST
***************************************

*.CALIBRE ABORT_INFO SOFTCHK
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lcesd1_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT lcesd2_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_shield PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_wos PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_x_40k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_x_40k PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_x_40k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nr36 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_w40 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT tsmc_c018_sealring_corner_1p6m
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT tsmc_c018_seal_ring_edge_1p6m
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=23093 EP=0 IP=93 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27
** N=11242 EP=0 IP=54 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=422 EP=0 IP=42 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=677 EP=0 IP=36 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=541 EP=0 IP=54 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=547 EP=0 IP=51 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=10106 EP=0 IP=54 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21
** N=23120 EP=0 IP=93 FDC=0
.ENDS
***************************************
.SUBCKT padbox
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pad_in VSS pad VDD DataIn
** N=24 EP=4 IP=1 FDC=96
M0 VSS VSS 7 VSS N L=3.5e-07 W=9e-06 $X=5700 $Y=147100 $D=0
M1 8 7 VSS VSS N L=3.5e-07 W=9e-06 $X=8100 $Y=147100 $D=0
M2 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=13200 $Y=147100 $D=0
M3 10 VSS VSS VSS N L=3.5e-07 W=9e-06 $X=15600 $Y=147100 $D=0
M4 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=191300 $D=0
M5 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=196210 $D=0
M6 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=197780 $D=0
M7 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=202690 $D=0
M8 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=204260 $D=0
M9 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=209170 $D=0
M10 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=210740 $D=0
M11 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=215650 $D=0
M12 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=217220 $D=0
M13 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=222130 $D=0
M14 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=18000 $Y=147100 $D=0
M15 10 VSS VSS VSS N L=3.5e-07 W=9e-06 $X=20400 $Y=147100 $D=0
M16 VSS VSS 10 VSS N L=3.5e-07 W=9e-06 $X=22800 $Y=147100 $D=0
M17 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=25200 $Y=147100 $D=0
M18 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=27600 $Y=147100 $D=0
M19 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=30000 $Y=147100 $D=0
M20 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=32400 $Y=147100 $D=0
M21 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=34800 $Y=147100 $D=0
M22 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=37200 $Y=147100 $D=0
M23 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=39600 $Y=147100 $D=0
M24 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=42000 $Y=147100 $D=0
M25 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=44400 $Y=147100 $D=0
M26 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=191300 $D=0
M27 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=196210 $D=0
M28 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=197780 $D=0
M29 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=202690 $D=0
M30 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=204260 $D=0
M31 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=209170 $D=0
M32 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=210740 $D=0
M33 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=215650 $D=0
M34 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=217220 $D=0
M35 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=222130 $D=0
M36 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=59400 $Y=146950 $D=0
M37 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=61800 $Y=146950 $D=0
M38 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=64200 $Y=146950 $D=0
M39 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=66600 $Y=146950 $D=0
M40 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=69000 $Y=146950 $D=0
M41 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=71400 $Y=146950 $D=0
M42 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=73800 $Y=146950 $D=0
M43 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=76200 $Y=146950 $D=0
M44 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=78600 $Y=146950 $D=0
M45 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=81000 $Y=146950 $D=0
M46 DataIn 11 VSS VSS N L=3.5e-07 W=9e-06 $X=83400 $Y=146950 $D=0
M47 VSS 11 DataIn VSS N L=3.5e-07 W=9e-06 $X=85800 $Y=146950 $D=0
M48 VDD VSS 7 VDD P L=3.5e-07 W=1.56e-05 $X=5700 $Y=165550 $D=16
M49 8 7 VDD VDD P L=3.5e-07 W=1.56e-05 $X=8100 $Y=165550 $D=16
M50 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=13200 $Y=165550 $D=16
M51 9 VSS VDD VDD P L=3.5e-07 W=1.56e-05 $X=15600 $Y=165550 $D=16
M52 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=97085 $D=16
M53 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=101995 $D=16
M54 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=103565 $D=16
M55 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=108475 $D=16
M56 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=110045 $D=16
M57 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=114955 $D=16
M58 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=116525 $D=16
M59 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=121435 $D=16
M60 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=123005 $D=16
M61 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=127915 $D=16
M62 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=18000 $Y=165550 $D=16
M63 9 VSS VDD VDD P L=3.5e-07 W=1.56e-05 $X=20400 $Y=165550 $D=16
M64 VDD VSS 9 VDD P L=3.5e-07 W=1.56e-05 $X=22800 $Y=165550 $D=16
M65 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=25200 $Y=165550 $D=16
M66 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=27600 $Y=165550 $D=16
M67 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=30000 $Y=165550 $D=16
M68 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=32400 $Y=165550 $D=16
M69 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=34800 $Y=165550 $D=16
M70 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=37200 $Y=165550 $D=16
M71 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=39600 $Y=165550 $D=16
M72 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=42000 $Y=165550 $D=16
M73 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=44400 $Y=165550 $D=16
M74 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=97085 $D=16
M75 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=101995 $D=16
M76 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=103565 $D=16
M77 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=108475 $D=16
M78 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=110045 $D=16
M79 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=114955 $D=16
M80 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=116525 $D=16
M81 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=121435 $D=16
M82 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=123005 $D=16
M83 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=127915 $D=16
M84 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=59400 $Y=165550 $D=16
M85 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=61800 $Y=165550 $D=16
M86 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=64200 $Y=165550 $D=16
M87 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=66600 $Y=165550 $D=16
M88 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=69000 $Y=165550 $D=16
M89 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=71400 $Y=165550 $D=16
M90 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=73800 $Y=165550 $D=16
M91 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=76200 $Y=165550 $D=16
M92 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=78600 $Y=165550 $D=16
M93 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=81000 $Y=165550 $D=16
M94 DataIn 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=83400 $Y=165550 $D=16
M95 VDD 11 DataIn VDD P L=3.5e-07 W=1.56e-05 $X=85800 $Y=165550 $D=16
.ENDS
***************************************
.SUBCKT pad_out VDD DataOut pad VSS
** N=25 EP=4 IP=1 FDC=96
M0 VSS VDD 7 VSS N L=3.5e-07 W=9e-06 $X=5700 $Y=147100 $D=0
M1 8 7 VSS VSS N L=3.5e-07 W=9e-06 $X=8100 $Y=147100 $D=0
M2 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=13200 $Y=147100 $D=0
M3 10 DataOut VSS VSS N L=3.5e-07 W=9e-06 $X=15600 $Y=147100 $D=0
M4 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=191300 $D=0
M5 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=196210 $D=0
M6 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=197780 $D=0
M7 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=202690 $D=0
M8 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=204260 $D=0
M9 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=209170 $D=0
M10 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=210740 $D=0
M11 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=215650 $D=0
M12 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=217220 $D=0
M13 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=15770 $Y=222130 $D=0
M14 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=18000 $Y=147100 $D=0
M15 10 DataOut VSS VSS N L=3.5e-07 W=9e-06 $X=20400 $Y=147100 $D=0
M16 VSS DataOut 10 VSS N L=3.5e-07 W=9e-06 $X=22800 $Y=147100 $D=0
M17 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=25200 $Y=147100 $D=0
M18 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=27600 $Y=147100 $D=0
M19 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=30000 $Y=147100 $D=0
M20 VSS 7 10 VSS N L=3.5e-07 W=9e-06 $X=32400 $Y=147100 $D=0
M21 10 7 VSS VSS N L=3.5e-07 W=9e-06 $X=34800 $Y=147100 $D=0
M22 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=37200 $Y=147100 $D=0
M23 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=39600 $Y=147100 $D=0
M24 9 8 10 VSS N L=3.5e-07 W=9e-06 $X=42000 $Y=147100 $D=0
M25 10 8 9 VSS N L=3.5e-07 W=9e-06 $X=44400 $Y=147100 $D=0
M26 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=191300 $D=0
M27 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=196210 $D=0
M28 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=197780 $D=0
M29 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=202690 $D=0
M30 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=204260 $D=0
M31 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=209170 $D=0
M32 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=210740 $D=0
M33 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=215650 $D=0
M34 pad 10 VSS VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=217220 $D=0
M35 VSS 10 pad VSS N L=3.5e-07 W=2e-05 $X=54230 $Y=222130 $D=0
M36 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=59400 $Y=146950 $D=0
M37 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=61800 $Y=146950 $D=0
M38 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=64200 $Y=146950 $D=0
M39 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=66600 $Y=146950 $D=0
M40 11 pad VSS VSS N L=3.5e-07 W=9e-06 $X=69000 $Y=146950 $D=0
M41 VSS pad 11 VSS N L=3.5e-07 W=9e-06 $X=71400 $Y=146950 $D=0
M42 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=73800 $Y=146950 $D=0
M43 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=76200 $Y=146950 $D=0
M44 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=78600 $Y=146950 $D=0
M45 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=81000 $Y=146950 $D=0
M46 12 11 VSS VSS N L=3.5e-07 W=9e-06 $X=83400 $Y=146950 $D=0
M47 VSS 11 12 VSS N L=3.5e-07 W=9e-06 $X=85800 $Y=146950 $D=0
M48 VDD VDD 7 VDD P L=3.5e-07 W=1.56e-05 $X=5700 $Y=165550 $D=16
M49 8 7 VDD VDD P L=3.5e-07 W=1.56e-05 $X=8100 $Y=165550 $D=16
M50 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=13200 $Y=165550 $D=16
M51 9 DataOut VDD VDD P L=3.5e-07 W=1.56e-05 $X=15600 $Y=165550 $D=16
M52 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=97085 $D=16
M53 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=101995 $D=16
M54 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=103565 $D=16
M55 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=108475 $D=16
M56 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=110045 $D=16
M57 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=114955 $D=16
M58 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=116525 $D=16
M59 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=121435 $D=16
M60 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=123005 $D=16
M61 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=15795 $Y=127915 $D=16
M62 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=18000 $Y=165550 $D=16
M63 9 DataOut VDD VDD P L=3.5e-07 W=1.56e-05 $X=20400 $Y=165550 $D=16
M64 VDD DataOut 9 VDD P L=3.5e-07 W=1.56e-05 $X=22800 $Y=165550 $D=16
M65 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=25200 $Y=165550 $D=16
M66 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=27600 $Y=165550 $D=16
M67 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=30000 $Y=165550 $D=16
M68 VDD 8 9 VDD P L=3.5e-07 W=1.56e-05 $X=32400 $Y=165550 $D=16
M69 9 8 VDD VDD P L=3.5e-07 W=1.56e-05 $X=34800 $Y=165550 $D=16
M70 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=37200 $Y=165550 $D=16
M71 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=39600 $Y=165550 $D=16
M72 10 7 9 VDD P L=3.5e-07 W=1.56e-05 $X=42000 $Y=165550 $D=16
M73 9 7 10 VDD P L=3.5e-07 W=1.56e-05 $X=44400 $Y=165550 $D=16
M74 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=97085 $D=16
M75 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=101995 $D=16
M76 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=103565 $D=16
M77 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=108475 $D=16
M78 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=110045 $D=16
M79 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=114955 $D=16
M80 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=116525 $D=16
M81 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=121435 $D=16
M82 pad 9 VDD VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=123005 $D=16
M83 VDD 9 pad VDD P L=3.5e-07 W=2e-05 $X=53330 $Y=127915 $D=16
M84 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=59400 $Y=165550 $D=16
M85 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=61800 $Y=165550 $D=16
M86 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=64200 $Y=165550 $D=16
M87 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=66600 $Y=165550 $D=16
M88 11 pad VDD VDD P L=3.5e-07 W=1.56e-05 $X=69000 $Y=165550 $D=16
M89 VDD pad 11 VDD P L=3.5e-07 W=1.56e-05 $X=71400 $Y=165550 $D=16
M90 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=73800 $Y=165550 $D=16
M91 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=76200 $Y=165550 $D=16
M92 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=78600 $Y=165550 $D=16
M93 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=81000 $Y=165550 $D=16
M94 12 11 VDD VDD P L=3.5e-07 W=1.56e-05 $X=83400 $Y=165550 $D=16
M95 VDD 11 12 VDD P L=3.5e-07 W=1.56e-05 $X=85800 $Y=165550 $D=16
.ENDS
***************************************
.SUBCKT ICV_95 33 34 35 165 166
** N=6814 EP=5 IP=12 FDC=192
X0 33 165 34 35 pad_in $T=0 323200 0 270 $X=0 $Y=232300
X1 34 33 166 33 pad_out $T=0 413200 0 270 $X=0 $Y=322300
.ENDS
***************************************
.SUBCKT ICV_34 22 23 24 110
** N=3216 EP=4 IP=6 FDC=96
X0 23 24 110 22 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_94
** N=171 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4 VSS VDD
** N=425 EP=2 IP=1 FDC=1
D0 VSS VDD pdio_m AREA=9e-10 PJ=0.00012 $X=8570 $Y=96300 $D=31
.ENDS
***************************************
.SUBCKT ICV_32 21 22 89
** N=3055 EP=3 IP=6 FDC=96
X0 22 21 89 21 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_93 25 26 114 115
** N=6552 EP=4 IP=12 FDC=192
X0 26 25 114 25 pad_out $T=0 773200 0 270 $X=0 $Y=682300
X1 26 25 115 25 pad_out $T=0 863200 0 270 $X=0 $Y=772300
.ENDS
***************************************
.SUBCKT ICV_92 33 34 143 144
** N=6272 EP=4 IP=12 FDC=192
X0 34 33 143 33 pad_out $T=0 953200 0 270 $X=0 $Y=862300
X1 34 33 144 33 pad_out $T=0 1043200 0 270 $X=0 $Y=952300
.ENDS
***************************************
.SUBCKT ICV_30 22 23 94
** N=2998 EP=3 IP=6 FDC=96
X0 23 22 94 22 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_91 24 25 112 113
** N=6588 EP=4 IP=12 FDC=192
X0 25 24 112 24 pad_out $T=0 1223200 0 270 $X=0 $Y=1132300
X1 25 24 113 24 pad_out $T=0 1313200 0 270 $X=0 $Y=1222300
.ENDS
***************************************
.SUBCKT pad_corner
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_90 11 18 261
** N=6826 EP=3 IP=10 FDC=96
X0 18 11 261 11 pad_out $T=0 1403200 0 270 $X=0 $Y=1312300
.ENDS
***************************************
.SUBCKT ICV_96
** N=3495 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35 224 254 255 332 363 1597 1598 1599 1600 1601 1602 1603 1604 1605 1606 1607 1608 1609 1610
** N=82969 EP=19 IP=88 FDC=1344
X0 224 1597 254 255 pad_in $T=323200 1636400 0 180 $X=232300 $Y=1402300
X1 254 224 1598 224 pad_out $T=503200 1636400 0 180 $X=412300 $Y=1402300
X2 254 224 1599 224 pad_out $T=593200 1636400 0 180 $X=502300 $Y=1402300
X3 254 224 1600 224 pad_out $T=683200 1636400 0 180 $X=592300 $Y=1402300
X4 254 332 1601 224 pad_out $T=773200 1636400 0 180 $X=682300 $Y=1402300
X5 254 224 1602 224 pad_out $T=863200 1636400 0 180 $X=772300 $Y=1402300
X6 254 363 1603 224 pad_out $T=953200 1636400 0 180 $X=862300 $Y=1402300
X7 254 224 1604 224 pad_out $T=1043200 1636400 0 180 $X=952300 $Y=1402300
X8 254 224 1605 224 pad_out $T=1133200 1636400 0 180 $X=1042300 $Y=1402300
X9 254 224 1606 224 pad_out $T=1223200 1636400 0 180 $X=1132300 $Y=1402300
X10 254 224 1607 224 pad_out $T=1313200 1636400 0 180 $X=1222300 $Y=1402300
X11 254 224 1608 224 pad_out $T=1403200 1636400 0 180 $X=1312300 $Y=1402300
X12 254 224 1609 224 pad_out $T=1493200 1636400 0 180 $X=1402300 $Y=1402300
X13 254 224 1610 224 pad_out $T=1726400 1313200 0 90 $X=1492300 $Y=1312300
.ENDS
***************************************
.SUBCKT pad_fill_4
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT pad_fill_01
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_88
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT pad_fill_005
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_86
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_87
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_89 22 55 56 60 87 95 927 928 929 930 931 932 933 934 935 936 937 938 939
** N=56150 EP=19 IP=418 FDC=1248
X0 22 927 55 56 pad_in $T=239630 0 0 0 $X=238730 $Y=0
X1 22 928 55 60 pad_in $T=336060 0 0 0 $X=335160 $Y=0
X2 22 929 55 87 pad_in $T=1011050 0 0 0 $X=1010150 $Y=0
X3 55 22 930 22 pad_out $T=432490 0 0 0 $X=431590 $Y=0
X4 55 22 931 22 pad_out $T=528920 0 0 0 $X=528020 $Y=0
X5 55 22 932 22 pad_out $T=625350 0 0 0 $X=624450 $Y=0
X6 55 22 933 22 pad_out $T=721775 0 0 0 $X=720875 $Y=0
X7 55 22 934 22 pad_out $T=818200 0 0 0 $X=817300 $Y=0
X8 55 22 935 22 pad_out $T=914625 0 0 0 $X=913725 $Y=0
X9 55 22 936 22 pad_out $T=1107480 0 0 0 $X=1106580 $Y=0
X10 55 95 937 22 pad_out $T=1203910 0 0 0 $X=1203010 $Y=0
X11 55 22 938 22 pad_out $T=1300340 0 0 0 $X=1299440 $Y=0
X12 55 22 939 22 pad_out $T=1396770 0 0 0 $X=1395870 $Y=0
.ENDS
***************************************
.SUBCKT FILL32
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_70
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_74
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_84
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_41
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_42
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_43
** N=5 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_44
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_83
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_58
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT FILL16
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL8
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_56
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_78
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT DFFQSRX1 D CLK SETB RESETB VSS VDD Q
** N=34 EP=7 IP=0 FDC=40
M0 VSS D 20 VSS N L=1.8e-07 W=2.2e-07 $X=945 $Y=750 $D=0
M1 10 CLK VSS VSS N L=1.8e-07 W=2.2e-07 $X=1745 $Y=750 $D=0
M2 11 10 20 VSS N L=1.8e-07 W=2.2e-07 $X=3245 $Y=755 $D=0
M3 12 11 VSS VSS N L=1.8e-07 W=2.2e-07 $X=4745 $Y=755 $D=0
M4 13 12 VSS VSS N L=1.8e-07 W=2.2e-07 $X=6250 $Y=760 $D=0
M5 VSS 14 13 VSS N L=1.8e-07 W=2.2e-07 $X=7050 $Y=760 $D=0
M6 15 13 VSS VSS N L=1.8e-07 W=2.2e-07 $X=7850 $Y=1120 $D=0
M7 VSS SETB 14 VSS N L=1.8e-07 W=2.2e-07 $X=9355 $Y=755 $D=0
M8 22 CLK 11 VSS N L=1.8e-07 W=2.2e-07 $X=10860 $Y=750 $D=0
M9 33 15 VSS VSS N L=1.8e-07 W=4.4e-07 $X=12320 $Y=965 $D=0
M10 22 RESETB 33 VSS N L=1.8e-07 W=4.4e-07 $X=13040 $Y=965 $D=0
M11 16 CLK 15 VSS N L=1.8e-07 W=2.2e-07 $X=14500 $Y=755 $D=0
M12 34 16 VSS VSS N L=1.8e-07 W=4.4e-07 $X=15960 $Y=740 $D=0
M13 17 RESETB 34 VSS N L=1.8e-07 W=4.4e-07 $X=16680 $Y=740 $D=0
M14 18 17 VSS VSS N L=1.8e-07 W=2.2e-07 $X=18140 $Y=755 $D=0
M15 19 18 VSS VSS N L=1.8e-07 W=2.2e-07 $X=19640 $Y=755 $D=0
M16 VSS 14 19 VSS N L=1.8e-07 W=2.2e-07 $X=20440 $Y=755 $D=0
M17 24 19 VSS VSS N L=1.8e-07 W=2.2e-07 $X=21240 $Y=755 $D=0
M18 16 10 24 VSS N L=1.8e-07 W=2.2e-07 $X=22740 $Y=755 $D=0
M19 Q 17 VSS VSS N L=1.8e-07 W=2.2e-07 $X=24240 $Y=755 $D=0
M20 VDD D 20 VDD P L=1.8e-07 W=4.4e-07 $X=945 $Y=2705 $D=16
M21 10 CLK VDD VDD P L=1.8e-07 W=4.4e-07 $X=1665 $Y=2705 $D=16
M22 11 CLK 20 VDD P L=1.8e-07 W=4.4e-07 $X=3245 $Y=2725 $D=16
M23 12 11 VDD VDD P L=1.8e-07 W=4.4e-07 $X=4745 $Y=2725 $D=16
M24 21 12 13 VDD P L=1.8e-07 W=8.8e-07 $X=6250 $Y=2300 $D=16
M25 VDD 14 21 VDD P L=1.8e-07 W=8.8e-07 $X=6970 $Y=2300 $D=16
M26 15 13 VDD VDD P L=1.8e-07 W=4.4e-07 $X=7730 $Y=2520 $D=16
M27 VDD SETB 14 VDD P L=1.8e-07 W=4.4e-07 $X=9355 $Y=2535 $D=16
M28 22 10 11 VDD P L=1.8e-07 W=4.4e-07 $X=10815 $Y=2505 $D=16
M29 22 15 VDD VDD P L=1.8e-07 W=4.4e-07 $X=12320 $Y=2505 $D=16
M30 VDD RESETB 22 VDD P L=1.8e-07 W=4.4e-07 $X=13040 $Y=2505 $D=16
M31 16 10 15 VDD P L=1.8e-07 W=4.4e-07 $X=14500 $Y=2505 $D=16
M32 17 16 VDD VDD P L=1.8e-07 W=4.4e-07 $X=15960 $Y=2665 $D=16
M33 VDD RESETB 17 VDD P L=1.8e-07 W=4.4e-07 $X=16680 $Y=2665 $D=16
M34 18 17 VDD VDD P L=1.8e-07 W=4.4e-07 $X=18140 $Y=2725 $D=16
M35 23 18 19 VDD P L=1.8e-07 W=8.8e-07 $X=19640 $Y=2285 $D=16
M36 VDD 14 23 VDD P L=1.8e-07 W=8.8e-07 $X=20360 $Y=2285 $D=16
M37 24 19 VDD VDD P L=1.8e-07 W=4.4e-07 $X=21120 $Y=2505 $D=16
M38 16 CLK 24 VDD P L=1.8e-07 W=4.4e-07 $X=22740 $Y=2505 $D=16
M39 Q 17 VDD VDD P L=1.8e-07 W=4.4e-07 $X=24200 $Y=2505 $D=16
.ENDS
***************************************
.SUBCKT FILL4
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL1
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILL2
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_54
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT XOR2X1 B A VDD VSS Z
** N=11 EP=5 IP=0 FDC=10
M0 VSS B 10 VSS N L=1.8e-07 W=4.4e-07 $X=630 $Y=985 $D=0
M1 8 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=1350 $Y=985 $D=0
M2 9 8 10 VSS N L=1.8e-07 W=4.4e-07 $X=3205 $Y=1000 $D=0
M3 B A 9 VSS N L=1.8e-07 W=4.4e-07 $X=3925 $Y=1000 $D=0
M4 Z 9 VSS VSS N L=1.8e-07 W=4.4e-07 $X=5345 $Y=1000 $D=0
M5 VDD B 10 VDD P L=1.8e-07 W=4.4e-07 $X=630 $Y=2435 $D=16
M6 8 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1350 $Y=2435 $D=16
M7 9 A 10 VDD P L=1.8e-07 W=4.4e-07 $X=3205 $Y=2435 $D=16
M8 B 8 9 VDD P L=1.8e-07 W=4.4e-07 $X=3925 $Y=2435 $D=16
M9 Z 9 VDD VDD P L=1.8e-07 W=4.4e-07 $X=5345 $Y=2435 $D=16
.ENDS
***************************************
.SUBCKT AND2X1 A B VSS VDD Z
** N=10 EP=5 IP=0 FDC=6
M0 10 A 8 VSS N L=1.8e-07 W=4.4e-07 $X=905 $Y=750 $D=0
M1 VSS B 10 VSS N L=1.8e-07 W=4.4e-07 $X=1625 $Y=750 $D=0
M2 Z 8 VSS VSS N L=1.8e-07 W=2.2e-07 $X=2385 $Y=860 $D=0
M3 8 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=905 $Y=2670 $D=16
M4 VDD B 8 VDD P L=1.8e-07 W=4.4e-07 $X=1625 $Y=2670 $D=16
M5 Z 8 VDD VDD P L=1.8e-07 W=4.4e-07 $X=2385 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT ICV_76
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT OR2X1 A B VSS VDD Z
** N=12 EP=5 IP=0 FDC=6
M0 8 A VSS VSS N L=1.8e-07 W=2.2e-07 $X=835 $Y=760 $D=0
M1 VSS B 8 VSS N L=1.8e-07 W=2.2e-07 $X=1635 $Y=760 $D=0
M2 Z 8 VSS VSS N L=1.8e-07 W=2.2e-07 $X=2435 $Y=760 $D=0
M3 9 A 8 VDD P L=1.8e-07 W=8.8e-07 $X=835 $Y=2300 $D=16
M4 VDD B 9 VDD P L=1.8e-07 W=8.8e-07 $X=1555 $Y=2300 $D=16
M5 Z 8 VDD VDD P L=1.8e-07 W=4.4e-07 $X=2315 $Y=2520 $D=16
.ENDS
***************************************
.SUBCKT NAND3X1 A B C VSS VDD Z
** N=10 EP=6 IP=0 FDC=6
M0 9 A VSS VSS N L=1.8e-07 W=6.6e-07 $X=1210 $Y=745 $D=0
M1 10 B 9 VSS N L=1.8e-07 W=6.6e-07 $X=1930 $Y=745 $D=0
M2 Z C 10 VSS N L=1.8e-07 W=6.6e-07 $X=2650 $Y=745 $D=0
M3 Z A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1210 $Y=2670 $D=16
M4 VDD B Z VDD P L=1.8e-07 W=4.4e-07 $X=1930 $Y=2670 $D=16
M5 Z C VDD VDD P L=1.8e-07 W=4.4e-07 $X=2650 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT NOR2X1 A B VSS VDD Z
** N=10 EP=5 IP=0 FDC=4
M0 Z A VSS VSS N L=1.8e-07 W=2.2e-07 $X=925 $Y=760 $D=0
M1 VSS B Z VSS N L=1.8e-07 W=2.2e-07 $X=1725 $Y=760 $D=0
M2 8 A VDD VDD P L=1.8e-07 W=8.8e-07 $X=925 $Y=2300 $D=16
M3 Z B 8 VDD P L=1.8e-07 W=8.8e-07 $X=1645 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT ICV_63
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT INVX2 A VSS VDD Z
** N=6 EP=4 IP=0 FDC=2
M0 Z A VSS VSS N L=1.8e-07 W=4.4e-07 $X=740 $Y=740 $D=0
M1 Z A VDD VDD P L=1.8e-07 W=8.8e-07 $X=740 $Y=2300 $D=16
.ENDS
***************************************
.SUBCKT ICV_77
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT NAND2X1 A B VSS VDD Z
** N=9 EP=5 IP=0 FDC=4
M0 9 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=985 $Y=745 $D=0
M1 Z B 9 VSS N L=1.8e-07 W=4.4e-07 $X=1705 $Y=745 $D=0
M2 Z A VDD VDD P L=1.8e-07 W=4.4e-07 $X=985 $Y=2670 $D=16
M3 VDD B Z VDD P L=1.8e-07 W=4.4e-07 $X=1705 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT ICV_59
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_60
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_61
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT DFFQX1 CLK Q VDD D VSS
** N=16 EP=5 IP=0 FDC=18
M0 8 CLK VSS VSS N L=1.8e-07 W=2.2e-07 $X=870 $Y=750 $D=0
M1 9 8 D VSS N L=1.8e-07 W=2.2e-07 $X=2370 $Y=750 $D=0
M2 VSS 9 10 VSS N L=1.8e-07 W=2.2e-07 $X=3960 $Y=750 $D=0
M3 12 10 VSS VSS N L=1.8e-07 W=2.2e-07 $X=5720 $Y=750 $D=0
M4 9 CLK 12 VSS N L=1.8e-07 W=2.2e-07 $X=6755 $Y=750 $D=0
M5 11 CLK 10 VSS N L=1.8e-07 W=2.2e-07 $X=8440 $Y=750 $D=0
M6 13 8 11 VSS N L=1.8e-07 W=2.2e-07 $X=9640 $Y=750 $D=0
M7 VSS Q 13 VSS N L=1.8e-07 W=2.2e-07 $X=10440 $Y=750 $D=0
M8 Q 11 VSS VSS N L=1.8e-07 W=2.2e-07 $X=11240 $Y=750 $D=0
M9 8 CLK VDD VDD P L=1.8e-07 W=4.4e-07 $X=870 $Y=2670 $D=16
M10 9 CLK D VDD P L=1.8e-07 W=4.4e-07 $X=2460 $Y=2670 $D=16
M11 VDD 9 10 VDD P L=1.8e-07 W=4.4e-07 $X=3960 $Y=2670 $D=16
M12 12 10 VDD VDD P L=1.8e-07 W=4.4e-07 $X=5460 $Y=2670 $D=16
M13 9 8 12 VDD P L=1.8e-07 W=4.4e-07 $X=6180 $Y=2670 $D=16
M14 11 8 10 VDD P L=1.8e-07 W=4.4e-07 $X=7980 $Y=2670 $D=16
M15 13 CLK 11 VDD P L=1.8e-07 W=4.4e-07 $X=9780 $Y=2670 $D=16
M16 VDD Q 13 VDD P L=1.8e-07 W=4.4e-07 $X=10500 $Y=2670 $D=16
M17 Q 11 VDD VDD P L=1.8e-07 W=4.4e-07 $X=11220 $Y=2670 $D=16
.ENDS
***************************************
.SUBCKT ICV_80
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MUX2X1 A S B VSS VDD Z
** N=16 EP=6 IP=0 FDC=12
M0 VSS S 9 VSS N L=1.8e-07 W=4.4e-07 $X=940 $Y=960 $D=0
M1 15 A VSS VSS N L=1.8e-07 W=4.4e-07 $X=1660 $Y=960 $D=0
M2 10 9 15 VSS N L=1.8e-07 W=4.4e-07 $X=2380 $Y=960 $D=0
M3 16 S 10 VSS N L=1.8e-07 W=4.4e-07 $X=3100 $Y=960 $D=0
M4 VSS B 16 VSS N L=1.8e-07 W=4.4e-07 $X=3920 $Y=740 $D=0
M5 Z 10 VSS VSS N L=1.8e-07 W=4.4e-07 $X=4640 $Y=740 $D=0
M6 VDD S 9 VDD P L=1.8e-07 W=4.4e-07 $X=940 $Y=2520 $D=16
M7 11 A VDD VDD P L=1.8e-07 W=4.4e-07 $X=1660 $Y=2520 $D=16
M8 10 S 11 VDD P L=1.8e-07 W=4.4e-07 $X=2380 $Y=2520 $D=16
M9 12 9 10 VDD P L=1.8e-07 W=4.4e-07 $X=3100 $Y=2520 $D=16
M10 VDD B 12 VDD P L=1.8e-07 W=4.4e-07 $X=3920 $Y=2735 $D=16
M11 Z 10 VDD VDD P L=1.8e-07 W=4.4e-07 $X=4640 $Y=2735 $D=16
.ENDS
***************************************
.SUBCKT ICV_79
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_81
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_82
** N=5 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_85 50 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71
+ 72 73 74 75 76 77 78 79 80 81 82 83 84 130 132 1174 1175
** N=161802 EP=37 IP=4747 FDC=3012
X0 50 1174 53 23183 pad_in $T=1726400 233200 0 90 $X=1492300 $Y=232300
X1 50 1175 53 22949 pad_in $T=1726400 323200 0 90 $X=1492300 $Y=322300
X249 18199 80 130 53 50 53 18262 DFFQSRX1 $T=613440 434800 0 0 $X=613010 $Y=434410
X250 18508 80 130 53 50 53 18468 DFFQSRX1 $T=620160 434800 1 0 $X=619730 $Y=430245
X251 19206 80 130 53 50 53 18754 DFFQSRX1 $T=667200 434800 1 180 $X=641570 $Y=434410
X252 19559 80 130 53 50 53 19112 DFFQSRX1 $T=678960 426960 0 180 $X=653330 $Y=422405
X253 19812 80 130 53 50 53 19222 DFFQSRX1 $T=682880 419120 0 180 $X=657250 $Y=414565
X254 19854 80 130 53 50 53 19223 DFFQSRX1 $T=682880 458320 0 180 $X=657250 $Y=453765
X255 20138 80 130 53 50 53 19909 DFFQSRX1 $T=689040 411280 0 0 $X=688610 $Y=410890
X256 20611 80 130 53 50 53 20194 DFFQSRX1 $T=692400 419120 1 0 $X=691970 $Y=414565
X257 20748 80 130 53 50 53 20228 DFFQSRX1 $T=722640 426960 1 180 $X=697010 $Y=426570
X258 20700 80 130 53 50 53 20305 DFFQSRX1 $T=723200 442640 0 180 $X=697570 $Y=438085
X259 21133 80 79 53 50 53 21245 DFFQSRX1 $T=715360 411280 1 0 $X=714930 $Y=406725
X260 21218 80 79 53 50 53 21309 DFFQSRX1 $T=715920 403440 1 0 $X=715490 $Y=398885
X261 21243 80 79 53 50 53 21346 DFFQSRX1 $T=720960 387760 0 0 $X=720530 $Y=387370
X262 21418 80 79 53 50 53 21456 DFFQSRX1 $T=721520 364240 0 0 $X=721090 $Y=363850
X263 21323 80 79 53 50 53 21380 DFFQSRX1 $T=721520 372080 0 0 $X=721090 $Y=371690
X264 21322 80 79 53 50 53 21485 DFFQSRX1 $T=722080 356400 1 0 $X=721650 $Y=351845
X265 21285 80 79 53 50 53 21381 DFFQSRX1 $T=722640 426960 1 0 $X=722210 $Y=422405
X266 21296 80 79 53 50 53 21386 DFFQSRX1 $T=723200 442640 0 0 $X=722770 $Y=442250
X267 21417 80 79 53 50 53 21507 DFFQSRX1 $T=723200 458320 1 0 $X=722770 $Y=453765
X268 21697 80 79 53 50 53 21319 DFFQSRX1 $T=758480 395600 0 180 $X=732850 $Y=391045
X269 21704 80 79 53 50 53 21763 DFFQSRX1 $T=742240 348560 1 0 $X=741810 $Y=344005
X270 21713 80 79 53 50 53 21828 DFFQSRX1 $T=742240 434800 1 0 $X=741810 $Y=430245
X271 21727 80 79 53 50 53 21784 DFFQSRX1 $T=742240 442640 1 0 $X=741810 $Y=438085
X272 22123 80 79 53 50 53 21783 DFFQSRX1 $T=779760 356400 0 180 $X=754130 $Y=351845
X273 22070 80 79 53 50 53 21809 DFFQSRX1 $T=780880 379920 0 180 $X=755250 $Y=375365
X274 22107 80 79 53 50 53 21825 DFFQSRX1 $T=781440 379920 1 180 $X=755810 $Y=379530
X275 22147 80 79 53 50 53 21880 DFFQSRX1 $T=783680 395600 1 180 $X=758050 $Y=395210
X276 22054 80 79 53 50 53 21933 DFFQSRX1 $T=787040 419120 1 180 $X=761410 $Y=418730
X277 22393 80 79 53 50 53 21962 DFFQSRX1 $T=792640 411280 1 180 $X=767010 $Y=410890
X278 22610 80 79 53 50 53 22720 DFFQSRX1 $T=772480 387760 1 0 $X=772050 $Y=383205
X279 22750 80 53 79 50 53 22775 DFFQSRX1 $T=772480 403440 0 0 $X=772050 $Y=403050
X280 22533 80 79 53 50 53 22183 DFFQSRX1 $T=797680 426960 1 180 $X=772050 $Y=426570
X281 22679 80 79 53 50 53 22185 DFFQSRX1 $T=797680 450480 0 180 $X=772050 $Y=445925
X282 132 80 79 53 50 53 73 DFFQSRX1 $T=797680 458320 0 180 $X=772050 $Y=453765
X484 18299 18262 53 50 18199 XOR2X1 $T=629120 442640 1 180 $X=622530 $Y=442250
X485 19065 18754 53 50 19206 XOR2X1 $T=651520 442640 1 0 $X=651090 $Y=438085
X486 18943 63 53 50 62 XOR2X1 $T=657680 450480 1 180 $X=651090 $Y=450090
X487 19414 19112 53 50 19559 XOR2X1 $T=663840 426960 0 0 $X=663410 $Y=426570
X488 19645 19222 53 50 19786 XOR2X1 $T=673920 426960 0 0 $X=673490 $Y=426570
X489 19977 19223 53 50 19836 XOR2X1 $T=685120 450480 0 180 $X=678530 $Y=445925
X490 19927 19909 53 50 20138 XOR2X1 $T=684000 426960 1 0 $X=683570 $Y=422405
X491 20474 20194 53 50 20611 XOR2X1 $T=700800 426960 1 0 $X=700370 $Y=422405
X492 20559 20228 53 50 20748 XOR2X1 $T=705840 434800 0 0 $X=705410 $Y=434410
X493 21202 21245 53 50 21133 XOR2X1 $T=731600 419120 0 180 $X=725010 $Y=414565
X494 21358 21346 53 50 21243 XOR2X1 $T=736080 387760 0 180 $X=729490 $Y=383205
X495 21394 21380 53 50 21283 XOR2X1 $T=737760 379920 1 180 $X=731170 $Y=379530
X496 21375 21381 53 50 21285 XOR2X1 $T=737760 419120 1 180 $X=731170 $Y=418730
X497 21406 21386 53 50 21296 XOR2X1 $T=738320 442640 0 180 $X=731730 $Y=438085
X498 21493 21507 53 50 21417 XOR2X1 $T=743920 450480 1 180 $X=737330 $Y=450090
X499 21424 21485 53 50 21345 XOR2X1 $T=745040 364240 0 180 $X=738450 $Y=359685
X500 21829 21763 53 50 21701 XOR2X1 $T=757360 364240 0 180 $X=750770 $Y=359685
X501 21756 21828 53 50 21713 XOR2X1 $T=757920 426960 0 180 $X=751330 $Y=422405
X502 21743 69 53 50 68 XOR2X1 $T=758480 458320 0 180 $X=751890 $Y=453765
X503 21932 21880 53 50 22035 XOR2X1 $T=760160 403440 0 0 $X=759730 $Y=403050
X504 21905 21783 53 50 22123 XOR2X1 $T=764080 356400 0 0 $X=763650 $Y=356010
X505 21998 21933 53 50 22036 XOR2X1 $T=765200 419120 1 0 $X=764770 $Y=414565
X506 22171 21962 53 50 22393 XOR2X1 $T=776400 403440 1 0 $X=775970 $Y=398885
X507 22411 22183 53 50 22533 XOR2X1 $T=782000 434800 0 0 $X=781570 $Y=434410
X508 22476 22185 53 50 22679 XOR2X1 $T=787600 442640 1 0 $X=787170 $Y=438085
X509 22124 22720 53 50 22610 XOR2X1 $T=796560 387760 1 180 $X=789970 $Y=387370
X510 22820 22775 53 50 22750 XOR2X1 $T=802160 395600 1 180 $X=795570 $Y=395210
X511 18299 18262 50 53 54 AND2X1 $T=627440 450480 0 180 $X=623650 $Y=445925
X512 54 55 50 53 56 AND2X1 $T=624080 458320 1 0 $X=623650 $Y=453765
X513 18657 18468 50 53 18299 AND2X1 $T=641440 442640 1 180 $X=637650 $Y=442250
X514 60 18751 50 53 18943 AND2X1 $T=645360 450480 0 0 $X=644930 $Y=450090
X515 18943 63 50 53 19065 AND2X1 $T=659360 450480 0 180 $X=655570 $Y=445925
X516 19645 19222 50 53 19414 AND2X1 $T=673360 426960 1 180 $X=669570 $Y=426570
X517 64 19786 50 53 19812 AND2X1 $T=675600 434800 1 0 $X=675170 $Y=430245
X518 64 19836 50 53 19854 AND2X1 $T=682880 450480 1 180 $X=679090 $Y=450090
X519 19927 19871 50 53 19645 AND2X1 $T=683440 434800 0 180 $X=679650 $Y=430245
X520 19927 19909 50 53 19977 AND2X1 $T=684560 434800 0 0 $X=684130 $Y=434410
X521 20228 20194 50 53 20163 AND2X1 $T=693520 426960 1 180 $X=689730 $Y=426570
X522 65 66 50 53 20364 AND2X1 $T=694640 450480 1 0 $X=694210 $Y=445925
X523 64 20470 50 53 67 AND2X1 $T=699680 458320 1 0 $X=699250 $Y=453765
X524 20364 20305 50 53 20559 AND2X1 $T=701920 450480 1 0 $X=701490 $Y=445925
X525 20559 20228 50 53 20474 AND2X1 $T=710320 426960 0 180 $X=706530 $Y=422405
X526 21371 21345 50 53 21322 AND2X1 $T=736640 364240 0 180 $X=732850 $Y=359685
X527 21371 21283 50 53 21323 AND2X1 $T=736640 372080 0 180 $X=732850 $Y=367525
X528 21202 21245 50 53 21375 AND2X1 $T=733280 411280 0 0 $X=732850 $Y=410890
X529 21284 21309 50 53 21202 AND2X1 $T=737200 403440 1 180 $X=733410 $Y=403050
X530 21358 21346 50 53 21394 AND2X1 $T=741120 387760 0 180 $X=737330 $Y=383205
X531 21406 21386 50 53 21493 AND2X1 $T=738880 442640 1 0 $X=738450 $Y=438085
X532 21497 21527 50 53 21404 AND2X1 $T=745600 372080 0 180 $X=741810 $Y=367525
X533 21581 21319 50 53 21284 AND2X1 $T=747280 403440 1 180 $X=743490 $Y=403050
X534 21245 21381 50 53 21590 AND2X1 $T=743920 419120 1 0 $X=743490 $Y=414565
X535 21371 21671 50 53 21697 AND2X1 $T=748400 403440 1 0 $X=747970 $Y=398885
X536 21371 21701 50 53 21704 AND2X1 $T=754560 356400 0 180 $X=750770 $Y=351845
X537 21797 21784 50 53 21743 AND2X1 $T=761840 450480 0 180 $X=758050 $Y=445925
X538 21905 21783 50 53 21829 AND2X1 $T=762960 356400 1 180 $X=759170 $Y=356010
X539 21743 69 50 53 70 AND2X1 $T=759600 458320 1 0 $X=759170 $Y=453765
X540 21756 21828 50 53 21998 AND2X1 $T=761280 426960 1 0 $X=760850 $Y=422405
X541 21756 21887 50 53 21932 AND2X1 $T=761840 419120 1 0 $X=761410 $Y=414565
X542 21825 21809 50 53 21905 AND2X1 $T=762960 372080 1 0 $X=762530 $Y=367525
X543 21371 22036 50 53 22054 AND2X1 $T=764080 411280 0 0 $X=763650 $Y=410890
X544 21371 22035 50 53 22147 AND2X1 $T=768000 403440 0 0 $X=767570 $Y=403050
X545 21932 21880 50 53 22171 AND2X1 $T=769120 403440 1 0 $X=768690 $Y=398885
X546 22411 22183 50 53 22476 AND2X1 $T=782560 442640 1 0 $X=782130 $Y=438085
X547 74 22352 50 53 22411 AND2X1 $T=783120 450480 0 0 $X=782690 $Y=450090
X548 79 22653 50 53 22726 AND2X1 $T=798240 364240 0 180 $X=794450 $Y=359685
X549 22839 22868 50 53 22705 AND2X1 $T=798800 332880 1 0 $X=798370 $Y=328325
X550 79 22935 50 53 22836 AND2X1 $T=805520 372080 0 180 $X=801730 $Y=367525
X551 23002 22968 50 53 22945 AND2X1 $T=807200 317200 1 180 $X=803410 $Y=316810
X552 23086 23054 50 53 23034 AND2X1 $T=810560 348560 0 180 $X=806770 $Y=344005
X553 79 23133 50 53 22973 AND2X1 $T=810000 372080 0 0 $X=809570 $Y=371690
X554 22775 23184 50 53 23212 AND2X1 $T=812240 387760 1 0 $X=811810 $Y=383205
X555 23309 23357 50 53 23324 AND2X1 $T=819520 387760 1 0 $X=819090 $Y=383205
X556 23143 23109 50 53 22839 AND2X1 $T=825120 340720 1 180 $X=821330 $Y=340330
X590 18262 18421 50 53 18437 OR2X1 $T=629120 442640 0 0 $X=628690 $Y=442250
X591 55 18437 50 53 58 OR2X1 $T=629680 458320 1 0 $X=629250 $Y=453765
X592 18468 18531 50 53 18421 OR2X1 $T=636400 450480 0 180 $X=632610 $Y=445925
X593 18754 18966 50 53 18531 OR2X1 $T=650960 442640 1 180 $X=647170 $Y=442250
X594 63 19317 50 53 18966 OR2X1 $T=659360 450480 1 0 $X=658930 $Y=445925
X595 19112 19437 50 53 19317 OR2X1 $T=667200 442640 0 180 $X=663410 $Y=438085
X596 20194 20265 50 53 20107 OR2X1 $T=695760 434800 1 180 $X=691970 $Y=434410
X597 21386 21447 50 53 21472 OR2X1 $T=737760 434800 1 0 $X=737330 $Y=430245
X598 21309 21467 50 53 21468 OR2X1 $T=738880 403440 0 0 $X=738450 $Y=403050
X599 21245 21468 50 53 21487 OR2X1 $T=738880 411280 0 0 $X=738450 $Y=410890
X600 21381 21487 50 53 21447 OR2X1 $T=743360 419120 1 180 $X=739570 $Y=418730
X601 21507 21472 50 53 21578 OR2X1 $T=743360 434800 0 0 $X=742930 $Y=434410
X602 21670 21456 50 53 21609 OR2X1 $T=750640 372080 1 180 $X=746850 $Y=371690
X603 21828 21578 50 53 21898 OR2X1 $T=762400 434800 1 180 $X=758610 $Y=434410
X604 21784 21898 50 53 21992 OR2X1 $T=766880 450480 0 180 $X=763090 $Y=445925
X605 69 21992 50 53 71 OR2X1 $T=766880 458320 0 180 $X=763090 $Y=453765
X606 21825 22041 50 53 21371 OR2X1 $T=768000 387760 1 180 $X=764210 $Y=387370
X607 21962 22060 50 53 22041 OR2X1 $T=769120 411280 0 180 $X=765330 $Y=406725
X608 22185 75 50 53 22263 OR2X1 $T=779200 434800 1 180 $X=775410 $Y=434410
X609 77 22945 50 53 22970 OR2X1 $T=802160 325040 1 0 $X=801730 $Y=320485
X610 23109 23080 50 53 22736 OR2X1 $T=811120 340720 1 180 $X=807330 $Y=340330
X611 23200 23161 50 53 23068 OR2X1 $T=815040 356400 0 180 $X=811250 $Y=351845
X612 23050 23184 50 53 23275 OR2X1 $T=815040 364240 0 0 $X=814610 $Y=363850
X613 23297 23109 50 53 23200 OR2X1 $T=818960 325040 0 180 $X=815170 $Y=320485
X614 23109 23161 50 53 23423 OR2X1 $T=821200 356400 1 0 $X=820770 $Y=351845
X615 23306 23398 50 53 23469 OR2X1 $T=823440 395600 1 0 $X=823010 $Y=391045
X616 23306 23425 50 53 23376 OR2X1 $T=826800 403440 1 180 $X=823010 $Y=403050
X617 23274 23469 50 53 23375 OR2X1 $T=824560 395600 0 0 $X=824130 $Y=395210
X618 57 18468 18262 50 53 18489 NAND3X1 $T=630240 450480 0 0 $X=629810 $Y=450090
X619 18691 18754 63 50 53 19013 NAND3X1 $T=652080 450480 1 0 $X=651650 $Y=445925
X620 19625 19112 19222 50 53 19576 NAND3X1 $T=672800 442640 0 180 $X=668450 $Y=438085
X621 19767 19222 19223 50 53 19437 NAND3X1 $T=677840 442640 0 180 $X=673490 $Y=438085
X622 20163 66 20305 50 53 19910 NAND3X1 $T=691840 442640 1 0 $X=691410 $Y=438085
X623 20393 20398 66 50 53 20265 NAND3X1 $T=700800 434800 1 180 $X=696450 $Y=434410
X624 21547 21319 21380 50 53 21467 NAND3X1 $T=745600 387760 0 180 $X=741250 $Y=383205
X625 21566 21380 21346 50 53 21546 NAND3X1 $T=746720 379920 1 180 $X=742370 $Y=379530
X626 21590 21319 21309 50 53 21582 NAND3X1 $T=748400 411280 0 180 $X=744050 $Y=406725
X627 21796 21763 21485 50 53 21670 NAND3X1 $T=756240 372080 0 180 $X=751890 $Y=367525
X628 21905 21783 21763 50 53 21497 NAND3X1 $T=760720 364240 1 180 $X=756370 $Y=363850
X629 21830 21962 21880 50 53 21810 NAND3X1 $T=760160 411280 1 0 $X=759730 $Y=406725
X630 72 21784 69 50 53 22068 NAND3X1 $T=769680 450480 1 180 $X=765330 $Y=450090
X631 22236 21880 21933 50 53 22060 NAND3X1 $T=775840 419120 0 180 $X=771490 $Y=414565
X632 22285 22185 22183 50 53 22184 NAND3X1 $T=776400 442640 0 0 $X=775970 $Y=442250
X633 22718 22781 22819 50 53 22799 NAND3X1 $T=795440 348560 1 0 $X=795010 $Y=344005
X634 23068 23034 22920 50 53 22905 NAND3X1 $T=810000 348560 1 180 $X=805650 $Y=348170
X635 23085 23050 22942 50 53 23002 NAND3X1 $T=810560 325040 1 180 $X=806210 $Y=324650
X636 22839 23080 22977 50 53 23054 NAND3X1 $T=811680 332880 1 180 $X=807330 $Y=332490
X637 23126 23109 23183 50 53 22790 NAND3X1 $T=810560 317200 1 0 $X=810130 $Y=312645
X638 23126 23109 23108 50 53 23086 NAND3X1 $T=814480 325040 0 180 $X=810130 $Y=320485
X639 23200 23050 23143 50 53 22819 NAND3X1 $T=816160 348560 0 180 $X=811810 $Y=344005
X640 23161 23260 23275 50 53 23278 NAND3X1 $T=815040 356400 0 0 $X=814610 $Y=356010
X641 23120 23143 23323 50 53 23260 NAND3X1 $T=816160 356400 1 0 $X=815730 $Y=351845
X642 23324 23293 23158 50 53 23185 NAND3X1 $T=820640 403440 1 180 $X=816290 $Y=403050
X643 23126 22942 23297 50 53 23374 NAND3X1 $T=818960 325040 1 0 $X=818530 $Y=320485
X644 23324 23350 23440 50 53 23425 NAND3X1 $T=821200 403440 1 0 $X=820770 $Y=398885
X645 23322 23199 23143 50 53 23453 NAND3X1 $T=822320 332880 1 0 $X=821890 $Y=328325
X646 22970 23374 23453 50 53 23475 NAND3X1 $T=823440 325040 1 0 $X=823010 $Y=320485
X647 23488 23423 23534 50 53 23551 NAND3X1 $T=826240 348560 0 0 $X=825810 $Y=348170
X648 18527 18299 50 53 18508 NOR2X1 $T=635280 442640 1 180 $X=632050 $Y=442250
X649 18468 18657 50 53 18527 NOR2X1 $T=640880 442640 0 180 $X=637650 $Y=438085
X650 59 18489 50 53 18691 NOR2X1 $T=641440 450480 1 180 $X=638210 $Y=450090
X651 18489 18834 50 53 60 NOR2X1 $T=643120 450480 1 0 $X=642690 $Y=445925
X652 19013 18834 50 53 61 NOR2X1 $T=651520 450480 1 180 $X=648290 $Y=450090
X653 19611 19576 50 53 18657 NOR2X1 $T=672240 450480 0 180 $X=669010 $Y=445925
X654 19881 19910 50 53 19625 NOR2X1 $T=680080 442640 1 0 $X=679650 $Y=438085
X655 19910 19611 50 53 19927 NOR2X1 $T=686240 442640 0 0 $X=685810 $Y=442250
X656 19909 20107 50 53 19767 NOR2X1 $T=686800 434800 1 0 $X=686370 $Y=430245
X657 66 65 50 53 20352 NOR2X1 $T=695200 458320 1 0 $X=694770 $Y=453765
X658 20352 20364 50 53 20470 NOR2X1 $T=699680 450480 0 0 $X=699250 $Y=450090
X659 20305 20364 50 53 20612 NOR2X1 $T=705280 450480 0 0 $X=704850 $Y=450090
X660 20612 20559 50 53 20700 NOR2X1 $T=708080 450480 1 0 $X=707650 $Y=445925
X661 21230 21202 50 53 21218 NOR2X1 $T=730480 403440 1 180 $X=727250 $Y=403050
X662 21309 21284 50 53 21230 NOR2X1 $T=733840 403440 1 180 $X=730610 $Y=403050
X663 21404 21424 50 53 21418 NOR2X1 $T=736640 356400 0 0 $X=736210 $Y=356010
X664 21474 21497 50 53 21358 NOR2X1 $T=740000 379920 0 0 $X=739570 $Y=379530
X665 21319 21581 50 53 21567 NOR2X1 $T=744480 403440 1 0 $X=744050 $Y=398885
X666 21527 21497 50 53 21424 NOR2X1 $T=747280 364240 1 0 $X=746850 $Y=359685
X667 21346 21609 50 53 21547 NOR2X1 $T=747280 387760 0 0 $X=746850 $Y=387370
X668 21497 21546 50 53 21581 NOR2X1 $T=751760 379920 1 180 $X=748530 $Y=379530
X669 21567 21284 50 53 21671 NOR2X1 $T=748960 403440 0 0 $X=748530 $Y=403050
X670 21714 21743 50 53 21727 NOR2X1 $T=751200 450480 1 0 $X=750770 $Y=445925
X671 21582 21751 50 53 21756 NOR2X1 $T=752320 411280 0 0 $X=751890 $Y=410890
X672 21751 21810 50 53 21797 NOR2X1 $T=754000 419120 1 0 $X=753570 $Y=414565
X673 21784 21797 50 53 21714 NOR2X1 $T=754000 450480 1 0 $X=753570 $Y=445925
X674 21844 21582 50 53 21830 NOR2X1 $T=757920 411280 0 180 $X=754690 $Y=406725
X675 21783 21809 50 53 21796 NOR2X1 $T=758480 372080 1 0 $X=758050 $Y=367525
X676 22083 21905 50 53 22070 NOR2X1 $T=769120 364240 1 180 $X=765890 $Y=363850
X677 21825 22124 50 53 22107 NOR2X1 $T=768000 387760 0 0 $X=767570 $Y=387370
X678 21809 21825 50 53 22083 NOR2X1 $T=771360 372080 0 180 $X=768130 $Y=367525
X679 22184 22078 50 53 21406 NOR2X1 $T=773600 442640 0 180 $X=770370 $Y=438085
X680 22068 22078 50 53 74 NOR2X1 $T=774720 450480 1 180 $X=771490 $Y=450090
X681 76 22068 50 53 22285 NOR2X1 $T=779200 450480 1 180 $X=775970 $Y=450090
X682 22183 22263 50 53 22236 NOR2X1 $T=782000 434800 1 180 $X=778770 $Y=434410
X683 22601 22734 50 53 22717 NOR2X1 $T=793760 325040 1 0 $X=793330 $Y=320485
X684 22705 22735 50 53 22718 NOR2X1 $T=793760 332880 1 0 $X=793330 $Y=328325
X685 22736 22762 50 53 22749 NOR2X1 $T=794880 340720 1 0 $X=794450 $Y=336165
X686 78 22790 50 53 22735 NOR2X1 $T=796000 317200 1 0 $X=795570 $Y=312645
X687 78 22734 50 53 22817 NOR2X1 $T=797680 317200 0 0 $X=797250 $Y=316810
X688 22835 22749 50 53 22781 NOR2X1 $T=800480 340720 0 180 $X=797250 $Y=336165
X689 22800 22837 50 53 22820 NOR2X1 $T=797680 395600 1 0 $X=797250 $Y=391045
X690 22717 22817 50 53 22762 NOR2X1 $T=798240 325040 0 0 $X=797810 $Y=324650
X691 22949 77 50 53 22919 NOR2X1 $T=804960 340720 1 180 $X=801730 $Y=340330
X692 22919 22736 50 53 22904 NOR2X1 $T=802160 348560 1 0 $X=801730 $Y=344005
X693 22934 22960 50 53 22835 NOR2X1 $T=802720 340720 1 0 $X=802290 $Y=336165
X694 22949 23200 50 53 23085 NOR2X1 $T=813360 332880 0 0 $X=812930 $Y=332490
X695 23050 23200 50 53 23202 NOR2X1 $T=813360 340720 1 0 $X=812930 $Y=336165
X696 23183 23109 50 53 23069 NOR2X1 $T=814480 317200 1 0 $X=814050 $Y=312645
X697 23143 23050 50 53 23126 NOR2X1 $T=818960 348560 0 180 $X=815730 $Y=344005
X698 22942 23322 50 53 23302 NOR2X1 $T=817840 332880 1 0 $X=817410 $Y=328325
X699 23202 23302 50 53 22960 NOR2X1 $T=817840 340720 1 0 $X=817410 $Y=336165
X700 82 22934 50 53 23306 NOR2X1 $T=820640 372080 1 180 $X=817410 $Y=371690
X701 23050 23319 50 53 23399 NOR2X1 $T=824560 332880 1 180 $X=821330 $Y=332490
X702 82 23050 50 53 23274 NOR2X1 $T=826240 372080 1 180 $X=823010 $Y=371690
X703 23399 23475 50 53 23488 NOR2X1 $T=826800 332880 0 0 $X=826370 $Y=332490
X734 59 50 53 18751 INVX2 $T=640880 458320 1 0 $X=640450 $Y=453765
X735 18657 50 53 18834 INVX2 $T=643680 442640 0 0 $X=643250 $Y=442250
X736 19881 50 53 19871 INVX2 $T=681760 426960 1 180 $X=679650 $Y=426570
X737 65 50 53 19611 INVX2 $T=689600 450480 0 180 $X=687490 $Y=445925
X738 20305 50 53 20393 INVX2 $T=697440 442640 0 0 $X=697010 $Y=442250
X739 20228 50 53 20398 INVX2 $T=702480 434800 1 180 $X=700370 $Y=434410
X740 21474 50 53 21566 INVX2 $T=747280 379920 0 180 $X=745170 $Y=375365
X741 21456 50 53 21527 INVX2 $T=748400 364240 0 0 $X=747970 $Y=363850
X742 21581 50 53 21751 INVX2 $T=752320 411280 1 0 $X=751890 $Y=406725
X743 21844 50 53 21887 INVX2 $T=757920 411280 0 0 $X=757490 $Y=410890
X744 21797 50 53 22078 INVX2 $T=766880 450480 1 0 $X=766450 $Y=445925
X745 21371 50 53 22124 INVX2 $T=770800 395600 1 0 $X=770370 $Y=391045
X746 76 50 53 22352 INVX2 $T=779200 450480 0 0 $X=778770 $Y=450090
X747 77 50 53 22601 INVX2 $T=789280 325040 1 0 $X=788850 $Y=320485
X748 22720 50 53 22837 INVX2 $T=800480 387760 0 0 $X=800050 $Y=387370
X749 78 50 53 22942 INVX2 $T=802720 317200 1 0 $X=802290 $Y=312645
X750 22736 50 53 23120 INVX2 $T=810000 348560 0 0 $X=809570 $Y=348170
X751 82 50 53 79 INVX2 $T=810560 387760 1 0 $X=810130 $Y=383205
X752 23050 50 53 23080 INVX2 $T=811680 332880 1 0 $X=811250 $Y=328325
X753 22949 50 53 22977 INVX2 $T=813360 332880 1 180 $X=811250 $Y=332490
X754 23109 50 53 23184 INVX2 $T=813920 372080 0 0 $X=813490 $Y=371690
X755 23274 50 53 23293 INVX2 $T=817280 395600 0 0 $X=816850 $Y=395210
X756 23302 50 53 23319 INVX2 $T=818400 332880 0 0 $X=817970 $Y=332490
X757 22934 50 53 23143 INVX2 $T=818960 348560 1 0 $X=818530 $Y=344005
X758 23069 50 53 23322 INVX2 $T=819520 317200 1 0 $X=819090 $Y=312645
X759 23183 50 53 23297 INVX2 $T=825120 317200 1 180 $X=823010 $Y=316810
X782 19909 19223 50 53 19881 NAND2X1 $T=682880 434800 1 180 $X=679650 $Y=434410
X783 21456 21485 50 53 21474 NAND2X1 $T=739440 372080 1 0 $X=739010 $Y=367525
X784 21828 21933 50 53 21844 NAND2X1 $T=759040 419120 0 0 $X=758610 $Y=418730
X785 22904 22934 50 53 22920 NAND2X1 $T=801600 348560 0 0 $X=801170 $Y=348170
X786 22942 77 50 53 22933 NAND2X1 $T=804960 325040 1 180 $X=801730 $Y=324650
X787 22933 22977 50 53 22868 NAND2X1 $T=803280 332880 1 0 $X=802850 $Y=328325
X788 22934 22977 50 53 22734 NAND2X1 $T=805520 340720 1 0 $X=805090 $Y=336165
X789 22817 23069 50 53 22968 NAND2X1 $T=807200 317200 0 0 $X=806770 $Y=316810
X790 81 82 50 53 23158 NAND2X1 $T=811680 411280 1 0 $X=811250 $Y=406725
X791 22942 23183 50 53 23108 NAND2X1 $T=812800 317200 0 0 $X=812370 $Y=316810
X792 23080 22942 50 53 23199 NAND2X1 $T=813360 332880 1 0 $X=812930 $Y=328325
X793 23212 79 50 53 23309 NAND2X1 $T=817840 387760 0 0 $X=817410 $Y=387370
X794 23274 23109 50 53 23350 NAND2X1 $T=819520 395600 1 0 $X=819090 $Y=391045
X795 23126 23323 50 53 23161 NAND2X1 $T=820080 348560 0 0 $X=819650 $Y=348170
X796 23306 23109 50 53 23357 NAND2X1 $T=820080 379920 0 0 $X=819650 $Y=379530
X797 22839 22949 50 53 23534 NAND2X1 $T=826800 348560 1 0 $X=826370 $Y=344005
X798 84 82 50 53 23440 NAND2X1 $T=831280 403440 0 180 $X=828050 $Y=398885
X826 80 22653 53 22799 50 DFFQX1 $T=803280 356400 0 180 $X=790530 $Y=351845
X827 80 22934 53 22836 50 DFFQX1 $T=797680 372080 0 0 $X=797250 $Y=371690
X828 80 23050 53 22726 50 DFFQX1 $T=800480 364240 1 0 $X=800050 $Y=359685
X829 80 23133 53 22905 50 DFFQX1 $T=800480 364240 0 0 $X=800050 $Y=363850
X830 80 23109 53 22973 50 DFFQX1 $T=803280 379920 0 0 $X=802850 $Y=379530
X831 80 22800 53 22989 50 DFFQX1 $T=815600 395600 1 180 $X=802850 $Y=395210
X832 80 81 53 23185 50 DFFQX1 $T=816160 411280 1 180 $X=803410 $Y=410890
X833 80 83 53 23375 50 DFFQX1 $T=820080 411280 1 0 $X=819650 $Y=406725
X834 80 84 53 23376 50 DFFQX1 $T=820080 419120 1 0 $X=819650 $Y=414565
X835 80 23323 53 23278 50 DFFQX1 $T=832960 356400 1 180 $X=820210 $Y=356010
X836 80 22935 53 23551 50 DFFQX1 $T=832960 364240 1 180 $X=820210 $Y=363850
X853 22720 82 22800 50 53 22989 MUX2X1 $T=811120 387760 1 180 $X=805090 $Y=387370
X854 83 79 23212 50 53 23398 MUX2X1 $T=828480 387760 0 180 $X=822450 $Y=383205
.ENDS
***************************************
.SUBCKT ICV_69
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_71
** N=5 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_72
** N=7 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT ICV_73
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_65
** N=4 EP=0 IP=16 FDC=0
.ENDS
***************************************
.SUBCKT ICV_66
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_67
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_68
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_64
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_62
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_75 67 68 69 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99
+ 100 101 102 103 104 173 174 176 180 183 187 1126
** N=166381 EP=32 IP=1889 FDC=1504
M0 67 1711 68 67 N L=1.8e-07 W=2.2e-07 $X=625400 $Y=482600 $D=0
M1 69 1711 68 69 P L=1.8e-07 W=4.4e-07 $X=625400 $Y=484555 $D=16
X2 69 67 1126 67 pad_out $T=1726400 503200 0 90 $X=1492300 $Y=502300
X90 17261 174 68 69 67 69 83 DFFQSRX1 $T=611760 466160 0 0 $X=611330 $Y=465770
X91 173 174 176 69 67 69 1711 DFFQSRX1 $T=612320 489680 0 0 $X=611890 $Y=489290
X92 17298 174 68 69 67 69 17454 DFFQSRX1 $T=612880 481840 1 0 $X=612450 $Y=477285
X93 18348 174 68 69 67 69 17884 DFFQSRX1 $T=664960 481840 1 180 $X=639330 $Y=481450
X94 180 174 68 69 67 69 91 DFFQSRX1 $T=640880 458320 0 0 $X=640450 $Y=457930
X95 18437 174 68 69 67 69 17805 DFFQSRX1 $T=666080 474000 0 180 $X=640450 $Y=469445
X96 18438 174 68 69 67 69 17967 DFFQSRX1 $T=667200 489680 0 180 $X=641570 $Y=485125
X97 18457 174 68 69 67 69 17968 DFFQSRX1 $T=667200 505360 0 180 $X=641570 $Y=500805
X98 19235 174 68 69 67 69 19325 DFFQSRX1 $T=657680 497520 0 0 $X=657250 $Y=497130
X99 19159 174 68 69 67 69 19152 DFFQSRX1 $T=666080 474000 1 0 $X=665650 $Y=469445
X100 19423 174 68 69 67 69 18836 DFFQSRX1 $T=693520 466160 1 180 $X=667890 $Y=465770
X101 183 174 68 69 67 69 94 DFFQSRX1 $T=689040 458320 0 0 $X=688610 $Y=457930
X102 19630 174 68 69 67 69 19574 DFFQSRX1 $T=689040 505360 0 0 $X=688610 $Y=504970
X103 20370 174 68 69 67 69 19899 DFFQSRX1 $T=724320 466160 1 180 $X=698690 $Y=465770
X104 20298 174 68 69 67 69 19879 DFFQSRX1 $T=724320 474000 1 180 $X=698690 $Y=473610
X105 20403 174 68 69 67 69 19916 DFFQSRX1 $T=725440 497520 1 180 $X=699810 $Y=497130
X106 20792 174 68 69 67 69 20010 DFFQSRX1 $T=739440 481840 0 180 $X=713810 $Y=477285
X107 20751 174 68 69 67 69 20916 DFFQSRX1 $T=715920 489680 1 0 $X=715490 $Y=485125
X108 187 174 176 69 67 69 97 DFFQSRX1 $T=743360 458320 0 0 $X=742930 $Y=457930
X109 21873 174 176 69 67 69 22028 DFFQSRX1 $T=745040 474000 0 0 $X=744610 $Y=473610
X110 21894 174 176 69 67 69 22045 DFFQSRX1 $T=746160 489680 1 0 $X=745730 $Y=485125
X111 22954 174 176 69 67 69 22422 DFFQSRX1 $T=797680 474000 1 180 $X=772050 $Y=473610
X112 22977 174 176 69 67 69 104 DFFQSRX1 $T=772480 489680 0 0 $X=772050 $Y=489290
X199 84 83 69 67 17261 XOR2X1 $T=628000 458320 1 180 $X=621410 $Y=457930
X200 85 17454 69 67 17298 XOR2X1 $T=629120 474000 0 180 $X=622530 $Y=469445
X201 18187 17884 69 67 18348 XOR2X1 $T=648160 474000 0 0 $X=647730 $Y=473610
X202 89 17805 69 67 18437 XOR2X1 $T=650960 466160 1 0 $X=650530 $Y=461605
X203 90 17967 69 67 18438 XOR2X1 $T=650960 497520 1 0 $X=650530 $Y=492965
X204 18283 17968 69 67 18457 XOR2X1 $T=651520 513200 1 0 $X=651090 $Y=508645
X205 19212 19152 69 67 19037 XOR2X1 $T=680080 481840 1 180 $X=673490 $Y=481450
X206 19252 18836 69 67 19423 XOR2X1 $T=679520 466160 1 0 $X=679090 $Y=461605
X207 19558 19325 69 67 19268 XOR2X1 $T=690160 497520 0 180 $X=683570 $Y=492965
X208 20101 19916 69 67 20261 XOR2X1 $T=704720 497520 1 0 $X=704290 $Y=492965
X209 19939 19899 69 67 20370 XOR2X1 $T=708080 481840 0 0 $X=707650 $Y=481450
X210 20540 20916 69 67 20751 XOR2X1 $T=731040 497520 0 180 $X=724450 $Y=492965
X211 22048 22028 69 67 21873 XOR2X1 $T=762400 466160 1 180 $X=755810 $Y=465770
X212 95 22045 69 67 21894 XOR2X1 $T=762960 481840 0 180 $X=756370 $Y=477285
X213 22101 21629 69 67 21874 XOR2X1 $T=764080 497520 0 180 $X=757490 $Y=492965
X214 22326 22349 69 67 22498 XOR2X1 $T=769120 505360 1 0 $X=768690 $Y=500805
X215 102 22422 69 67 22954 XOR2X1 $T=782560 466160 0 0 $X=782130 $Y=465770
X216 22857 100 69 67 103 XOR2X1 $T=788160 466160 1 0 $X=787730 $Y=461605
X217 83 17454 67 69 86 AND2X1 $T=633600 458320 1 180 $X=629810 $Y=457930
X218 89 17805 67 69 18187 AND2X1 $T=645920 466160 1 0 $X=645490 $Y=461605
X219 90 17967 67 69 18283 AND2X1 $T=654880 497520 1 180 $X=651090 $Y=497130
X220 92 19037 67 69 19159 AND2X1 $T=680640 481840 0 180 $X=676850 $Y=477285
X221 92 19268 67 69 19235 AND2X1 $T=682880 497520 0 180 $X=679090 $Y=492965
X222 19252 18836 67 69 19212 AND2X1 $T=683440 481840 1 180 $X=679650 $Y=481450
X223 19593 19597 67 69 19650 AND2X1 $T=694640 497520 1 0 $X=694210 $Y=492965
X224 20010 19879 67 69 19939 AND2X1 $T=703600 481840 0 180 $X=699810 $Y=477285
X225 19939 19899 67 69 20101 AND2X1 $T=709200 489680 0 180 $X=705410 $Y=485125
X226 92 20261 67 69 20403 AND2X1 $T=712000 497520 1 0 $X=711570 $Y=492965
X227 95 22045 67 69 22048 AND2X1 $T=762960 481840 1 0 $X=762530 $Y=477285
X228 22045 22028 67 69 98 AND2X1 $T=765760 466160 1 0 $X=765330 $Y=461605
X229 102 22422 67 69 22857 AND2X1 $T=782560 466160 1 0 $X=782130 $Y=461605
X230 17454 87 67 69 17644 OR2X1 $T=630240 474000 1 0 $X=629810 $Y=469445
X231 17805 17644 67 69 17902 OR2X1 $T=637520 474000 1 0 $X=637090 $Y=469445
X232 17884 17902 67 69 18111 OR2X1 $T=643680 474000 0 0 $X=643250 $Y=473610
X233 20010 19133 67 69 92 OR2X1 $T=703040 497520 0 180 $X=699250 $Y=492965
X234 22028 96 67 69 22209 OR2X1 $T=763520 466160 0 0 $X=763090 $Y=465770
X235 22045 22209 67 69 22397 OR2X1 $T=769120 466160 0 0 $X=768690 $Y=465770
X236 22349 22250 67 69 22494 OR2X1 $T=771920 497520 1 0 $X=771490 $Y=492965
X237 100 22487 67 69 99 OR2X1 $T=777520 458320 1 180 $X=773730 $Y=457930
X238 22422 22397 67 69 22487 OR2X1 $T=777520 466160 0 180 $X=773730 $Y=461605
X239 18496 19106 19152 67 69 19133 NAND3X1 $T=673920 497520 1 0 $X=673490 $Y=492965
X240 19400 19152 18836 67 69 19362 NAND3X1 $T=685680 481840 0 180 $X=681330 $Y=477285
X241 19824 19871 19916 67 69 19745 NAND3X1 $T=696320 481840 0 0 $X=695890 $Y=481450
X242 19939 19899 19916 67 69 19593 NAND3X1 $T=704720 489680 0 180 $X=700370 $Y=485125
X243 17967 17968 67 69 18496 NOR2X1 $T=657120 497520 1 0 $X=656690 $Y=492965
X244 18836 19229 67 69 19106 NOR2X1 $T=677840 489680 1 0 $X=677410 $Y=485125
X245 19593 19362 67 69 93 NOR2X1 $T=691280 481840 0 180 $X=688050 $Y=477285
X246 19469 19593 67 69 19252 NOR2X1 $T=688480 481840 0 0 $X=688050 $Y=481450
X247 19650 19558 67 69 19630 NOR2X1 $T=692960 497520 0 180 $X=689730 $Y=492965
X248 19574 19745 67 69 19363 NOR2X1 $T=692960 489680 1 0 $X=692530 $Y=485125
X249 19597 19593 67 69 19558 NOR2X1 $T=695200 489680 0 0 $X=694770 $Y=489290
X250 19879 18111 67 69 19824 NOR2X1 $T=699680 481840 0 180 $X=696450 $Y=477285
X251 19879 20010 67 69 20152 NOR2X1 $T=705840 481840 1 0 $X=705410 $Y=477285
X252 20152 19939 67 69 20298 NOR2X1 $T=709760 481840 1 0 $X=709330 $Y=477285
X253 20010 20540 67 69 20792 NOR2X1 $T=724880 481840 0 0 $X=724450 $Y=481450
X258 19469 67 69 19400 INVX2 $T=686240 481840 0 0 $X=685810 $Y=481450
X259 19574 67 69 19597 INVX2 $T=691840 489680 1 180 $X=689730 $Y=489290
X260 19899 67 69 19871 INVX2 $T=704720 481840 1 180 $X=702610 $Y=481450
X261 92 67 69 20540 INVX2 $T=717600 497520 1 0 $X=717170 $Y=492965
X262 20916 67 69 21212 INVX2 $T=736640 497520 1 0 $X=736210 $Y=492965
X263 21629 67 69 21465 INVX2 $T=750080 489680 1 180 $X=747970 $Y=489290
X264 22250 67 69 22326 INVX2 $T=772480 497520 1 180 $X=770370 $Y=497130
X265 17805 17884 67 69 88 NAND2X1 $T=641440 466160 1 0 $X=641010 $Y=461605
X266 19363 19325 67 69 19229 NAND2X1 $T=682880 489680 1 0 $X=682450 $Y=485125
X267 19574 19325 67 69 19469 NAND2X1 $T=690720 489680 0 180 $X=687490 $Y=485125
X268 22101 21629 67 69 22250 NAND2X1 $T=769120 497520 0 180 $X=765890 $Y=492965
X269 22422 100 67 69 101 NAND2X1 $T=777520 466160 1 0 $X=777090 $Y=461605
X277 21212 21629 69 21465 67 DFFQX1 $T=742800 497520 0 0 $X=742370 $Y=497130
X278 21212 22101 69 21874 67 DFFQX1 $T=754560 505360 1 0 $X=754130 $Y=500805
X279 21212 22349 69 22498 67 DFFQX1 $T=776400 505360 1 0 $X=775970 $Y=500805
X280 21212 22977 69 22494 67 DFFQX1 $T=778080 497520 0 0 $X=777650 $Y=497130
.ENDS
***************************************
.SUBCKT ICV_45
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_46
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_47
** N=7 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_48
** N=11 EP=0 IP=14 FDC=0
.ENDS
***************************************
.SUBCKT ICV_49
** N=19 EP=0 IP=22 FDC=0
.ENDS
***************************************
.SUBCKT ICV_50
** N=35 EP=0 IP=38 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36
** N=5 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37
** N=7 EP=0 IP=10 FDC=0
.ENDS
***************************************
.SUBCKT ICV_53 58 82 172 982 983
** N=165619 EP=5 IP=1047 FDC=192
X0 82 58 982 58 pad_out $T=1726400 683200 0 90 $X=1492300 $Y=682300
X1 82 172 983 58 pad_out $T=1726400 773200 0 90 $X=1492300 $Y=772300
.ENDS
***************************************
.SUBCKT ICV_52 49 71 207 974 975
** N=163766 EP=5 IP=1047 FDC=192
X0 71 49 974 49 pad_out $T=1726400 863200 0 90 $X=1492300 $Y=862300
X1 71 207 975 49 pad_out $T=1726400 953200 0 90 $X=1492300 $Y=952300
.ENDS
***************************************
.SUBCKT ICV_51 50 63 1536 1537
** N=198468 EP=4 IP=1506 FDC=192
X0 63 50 1536 50 pad_out $T=1726400 1133200 0 90 $X=1492300 $Y=1132300
X1 63 50 1537 50 pad_out $T=1726400 1223200 0 90 $X=1492300 $Y=1222300
.ENDS
***************************************
.SUBCKT ICV_5 VSS VDD
** N=506 EP=2 IP=1 FDC=1
D0 VSS VDD ndio_m AREA=9e-10 PJ=0.00012 $X=10780 $Y=193610 $D=30
.ENDS
***************************************
.SUBCKT ICV_33 22 23 129
** N=3361 EP=3 IP=6 FDC=96
X0 23 22 129 22 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_31 21 22 23 131
** N=3340 EP=4 IP=6 FDC=96
X0 22 23 131 21 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_29 22 23 127
** N=3328 EP=3 IP=6 FDC=96
X0 23 22 127 22 pad_out $T=0 0 0 0 $X=-900 $Y=0
.ENDS
***************************************
.SUBCKT ICV_1 VSS
** N=6528 EP=1 IP=11113 FDC=9126
X0 VSS VDD 2798 clk h0_4 ICV_95 $T=0 0 0 0 $X=0 $Y=232300
X1 VSS VDD 2328 h0_0 ICV_34 $T=0 503200 0 270 $X=0 $Y=412300
X3 VSS VDD ICV_4 $T=0 593200 0 270 $X=0 $Y=502300
X4 VSS VDD h1_5 ICV_32 $T=0 683200 0 270 $X=0 $Y=592300
X5 VSS VDD h1_1 m0_5 ICV_93 $T=0 0 0 0 $X=0 $Y=680200
X6 VSS VDD m0_1 m1_6 ICV_92 $T=0 0 0 0 $X=0 $Y=862300
X7 VSS VDD m1_2 ICV_30 $T=0 1133200 0 270 $X=0 $Y=1042300
X8 VSS VDD s0_6 s0_2 ICV_91 $T=0 0 0 0 $X=0 $Y=1130200
X9 VSS VDD s1_3 ICV_90 $T=0 0 0 0 $X=0 $Y=1312300
X11 VSS VDD 2310 2328 2357 btn_light h0_3 colon h1_4 h1_0 m0_4 m0_0 m1_5 m1_1 s0_5 s0_1 s1_6 s1_2 s1_5 ICV_35 $T=0 0 0 0 $X=232300 $Y=1312300
X12 VSS VDD 2440 2441 2453 2457 btn_mode btn_dec reset h0_5 h0_1 h1_6 h1_2 m0_6 m0_2 m1_3 s1_0 s0_3 s1_4 ICV_89 $T=0 0 0 0 $X=232600 $Y=0
X13 VSS VDD 2493 2494 2495 2496 2497 2498 2499 4235 3267 3268 4237 4238 2500 3270 3273 2501 3274 3275
+ 2502 2503 4247 4245 4246 2441 2440 4242 2798 2328 2453 2457 2357 4236 2504 btn_set btn_inc
+ ICV_85 $T=0 0 0 0 $X=234100 $Y=232300
X14 VSS 4236 VDD 2494 2493 2495 2496 2497 2498 2499 4235 3268 4237 4238 2500 3274 3275 2501 2502 4245
+ 2503 4246 4247 2504 3445 2310 2798 4242 3267 3270 3273 h0_2
+ ICV_75 $T=0 0 0 0 $X=234100 $Y=457930
X15 VSS VDD 2357 h1_3 m1_0 ICV_53 $T=0 0 0 0 $X=234100 $Y=665400
X16 VSS VDD 2457 m0_3 s0_0 ICV_52 $T=0 0 0 0 $X=234100 $Y=862300
X17 VSS VDD s1_1 s0_4 ICV_51 $T=0 0 0 0 $X=234100 $Y=1073125
X18 VSS VDD ICV_5 $T=413200 1636400 0 180 $X=322300 $Y=1402300
X19 VSS VDD h0_6 ICV_33 $T=1726400 413200 0 90 $X=1492300 $Y=412300
X20 VSS VDD 3445 light ICV_31 $T=1726400 593200 0 90 $X=1492300 $Y=592300
X21 VSS VDD m1_4 ICV_29 $T=1726400 1043200 0 90 $X=1492300 $Y=1042300
.ENDS
***************************************
.SUBCKT ICV_2
** N=2764 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=2630 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20
** N=85952 EP=0 IP=93 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=84431 EP=0 IP=93 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19
** N=13895 EP=0 IP=54 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=13159 EP=0 IP=54 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18
** N=6233 EP=0 IP=42 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17
** N=9780 EP=0 IP=36 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=7962 EP=0 IP=54 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=7997 EP=0 IP=51 FDC=0
.ENDS
***************************************
.SUBCKT sealring_merged
** N=3694 EP=0 IP=7445 FDC=9126
X8 738 ICV_1 $T=67345 198305 0 0 $X=67345 $Y=198305
*.CALIBRE WARNING SCONNECT SCONNECT conflict(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
